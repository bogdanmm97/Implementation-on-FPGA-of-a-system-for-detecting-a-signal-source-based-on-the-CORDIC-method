module conv_dec_ascii(
	input [16:0] d_in,
	input clk,
	input en_conv,
	input again,
	
	output en_crc,
	output [47:0] d_out
    );
	reg [23:0] reg_d_out_i = 24'b0;
	reg [23:0] reg_data_out_q = 24'b0;
	reg reg_en_crc = 1'b0;
	
	assign d_out = {reg_d_out_i,reg_data_out_q};
	assign en_crc = reg_en_crc;
	
	always @(posedge clk) begin
		if(en_conv) begin
			reg_en_crc <= 1'b1;
			case (d_in[16:10])
				7'd0: reg_d_out_i <= {3{8'b00110000}};
				7'd1: reg_d_out_i <= {{2{8'b00110000}},8'b00110001};					
				7'd2: reg_d_out_i <= {{2{8'b00110000}},8'b00110010};
				7'd3: reg_d_out_i<= {{2{8'b00110000}},8'b00110011};
				7'd4: reg_d_out_i <= {{2{8'b00110000}},8'b00110100};
				7'd5: reg_d_out_i <= {{2{8'b00110000}},8'b00110101};
				7'd6: reg_d_out_i <= {{2{8'b00110000}},8'b00110110};
				7'd7: reg_d_out_i  <= {{2{8'b00110000}},8'b00110111};
				7'd8: reg_d_out_i  <= {{2{8'b00110000}},8'b00111001};
				7'd9: reg_d_out_i  <= {{2{8'b00110000}},8'b00111001};
				7'd10: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110000};
				7'd11: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110001};
				7'd12: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110010};
				7'd13: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110011};
				7'd14: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110100};
				7'd15: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110101};
				7'd16: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110110};
				7'd17: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110111};
				7'd18: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00111000};
				7'd19: reg_d_out_i  <= {8'b00110000,8'b00110001,8'b00110001};
				7'd20: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110000};
				7'd21: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110001};
				7'd22: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110010};
				7'd23: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110011};
				7'd24: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110100};
				7'd25: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110101};
				7'd26: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110110};
				7'd27: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00110111};
				7'd28: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00111000};
				7'd29: reg_d_out_i  <= {8'b00110000,8'b00110010,8'b00111001};
				7'd30: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110000};
				7'd31: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110001};
				7'd32: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110010};
				7'd33: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110011};
				7'd34: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110100};
				7'd35: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110101};
				7'd36: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110110};
				7'd37: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00110111};
				7'd38: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00111000};
				7'd39: reg_d_out_i  <= {8'b00110000,8'b00110011,8'b00111001};
				7'd40: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110000};
				7'd41: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110001};
				7'd42: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110010};
				7'd43: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110011};
				7'd44: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110100};
				7'd45: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110101};
				7'd46: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110110};
				7'd47: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00110111};
				7'd48: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00111000};
				7'd49: reg_d_out_i  <= {8'b00110000,8'b00110100,8'b00111001};
				7'd50: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110000};
				7'd51: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110001};
				7'd52: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110010};
				7'd53: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110011};
				7'd54: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110100};
				7'd55: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110101};
				7'd56: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110110};
				7'd57: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00110111};
				7'd58: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00111000};
				7'd59: reg_d_out_i  <= {8'b00110000,8'b00110101,8'b00111001};
				7'd60: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110000};
				7'd61: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110001};
				7'd62: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110010};
				7'd63: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110011};
				7'd64: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110100};
				7'd65: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110101};
				7'd66: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110110};
				7'd67: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00110111};
				7'd68: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00111000};
				7'd69: reg_d_out_i  <= {8'b00110000,8'b00110110,8'b00111001};
				7'd70: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110000};
				7'd71: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110001};
				7'd72: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110010};
				7'd73: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110011};
				7'd74: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110100};
				7'd75: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110101};
				7'd76: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110110};
				7'd77: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00110111};
				7'd78: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00111000};
				7'd79: reg_d_out_i  <= {8'b00110000,8'b00110111,8'b00111001};
				7'd80: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110000};
				7'd81: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110001};
				7'd82: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110010};
				7'd83: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110011};
				7'd84: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110100};
				7'd85: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110101};
				7'd86: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110110};
				7'd87: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00110111};
				7'd88: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00111000};
				7'd89: reg_d_out_i  <= {8'b00110000,8'b00111000,8'b00111001};
				7'd90: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110000};
				7'd91: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110001};
				7'd92: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110010};
				7'd93: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110011};
				7'd94: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110100};
				7'd95: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110110};
				7'd97: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00110111};
				7'd98: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00111000};
				7'd99: reg_d_out_i  <= {8'b00110000,8'b00111001,8'b00111001};
				7'd100: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110000};
				7'd101: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110001};
				7'd102: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110010};
				7'd103: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110011};
				7'd104: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110100};
				7'd105: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110101};
				7'd106: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110110};
				7'd107: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00110111};
				7'd108: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00111000};
				7'd109: reg_d_out_i  <= {8'b00110001,8'b00110000,8'b00111001};
				7'd110: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110000};
				7'd111: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110001};
				7'd112: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110010};
				7'd113: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110011};
				7'd114: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110100};
				7'd115: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110101};
				7'd116: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110110};
				7'd117: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00110111};
				7'd118: reg_d_out_i  <= {8'b00110001,8'b00110001,8'b00111001};
				7'd120: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110000};
				7'd121: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110001};
				7'd122: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110010};
				7'd123: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110011};
				7'd124: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110100};
				7'd125: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110101};
				7'd126: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110110};
				7'd127: reg_d_out_i  <= {8'b00110001,8'b00110010,8'b00110111};
			endcase
			case (d_in[9:0])
				  10'd000: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110000};
				  10'd001: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110001};
				  10'd002: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110010};
				  10'd003: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110011};
				  10'd004: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110100};
				  10'd005: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110101};
				  10'd006: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110110};
				  10'd007: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00110111};
				  10'd008: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00111000};
				  10'd009: reg_data_out_q <= {8'b00110000,8'b00110000,8'b00111001};
				  10'd010: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110000};
				  10'd011: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110001};
				  10'd012: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110010};
				  10'd013: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110011};
				  10'd014: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110100};
				  10'd015: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110101};
				  10'd016: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110110};
				  10'd017: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00110111};
				  10'd018: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00111000};
				  10'd019: reg_data_out_q <= {8'b00110000,8'b00110001,8'b00111001};
				  10'd020: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110000};
				  10'd021: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110001};
				  10'd022: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110010};
				  10'd023: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110011};
				  10'd024: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110100};
				  10'd025: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110101};
				  10'd026: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110110};
				  10'd027: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00110111};
				  10'd028: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00111000};
				  10'd029: reg_data_out_q <= {8'b00110000,8'b00110010,8'b00111001};
				  10'd030: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110000};
				  10'd031: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110001};
				  10'd032: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110010};
				  10'd033: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110011};
				  10'd034: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110100};
				  10'd035: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110101};
				  10'd036: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110110};
				  10'd037: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00110111};
				  10'd038: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00111000};
				  10'd039: reg_data_out_q <= {8'b00110000,8'b00110011,8'b00111001};
				  10'd040: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110000};
				  10'd041: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110001};
				  10'd041: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110001};
				  10'd042: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110010};
				  10'd043: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110011};
				  10'd044: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110100};
				  10'd045: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110101};
				  10'd046: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110110};
				  10'd047: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00110111};
				  10'd048: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00111000};
				  10'd049: reg_data_out_q <= {8'b00110000,8'b00110100,8'b00111001};
				  10'd050: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110000};
				  10'd051: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110001};
				  10'd052: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110010};
				  10'd053: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110011};
				  10'd054: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110100};
				  10'd055: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110101};
				  10'd056: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110110};
				  10'd057: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00110111};
				  10'd058: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00111000};
				  10'd059: reg_data_out_q <= {8'b00110000,8'b00110101,8'b00111001};
				  10'd060: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110000};
				  10'd061: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110001};
				  10'd062: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110010};
				  10'd063: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110011};
				  10'd064: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110100};
				  10'd065: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110101};
				  10'd066: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110110};
				  10'd067: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00110111};
				  10'd068: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00111000};
				  10'd069: reg_data_out_q <= {8'b00110000,8'b00110110,8'b00111001};
				  10'd070: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110000};
				  10'd071: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110001};
				  10'd072: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110010};
				  10'd073: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110011};
				  10'd074: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110100};
				  10'd075: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110101};
				  10'd076: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110110};
				  10'd077: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00110111};
				  10'd078: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00111000};
				  10'd079: reg_data_out_q <= {8'b00110000,8'b00110111,8'b00111001};
				  10'd080: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110000};
				  10'd081: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110001};
				  10'd082: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110010};
				  10'd083: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110011};
				  10'd083: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110011};
				  10'd084: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110100};
				  10'd085: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110101};
				  10'd086: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110110};
				  10'd087: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00110111};
				  10'd088: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00111000};
				  10'd089: reg_data_out_q <= {8'b00110000,8'b00111000,8'b00111001};
				  10'd090: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110000};
				  10'd091: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110001};
				  10'd092: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110010};
				  10'd093: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110011};
				  10'd094: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110100};
				  10'd095: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110101};
				  10'd096: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110110};
				  10'd097: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00110111};
				  10'd098: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00111000};
				  10'd099: reg_data_out_q <= {8'b00110000,8'b00111001,8'b00111001};
				  10'd100: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110000};
				  10'd101: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110001};
				  10'd102: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110010};
				  10'd103: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110011};
				  10'd104: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110100};
				  10'd105: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110101};
				  10'd106: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110110};
				  10'd107: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00110111};
				  10'd108: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00111000};
				  10'd109: reg_data_out_q <= {8'b00110001,8'b00110000,8'b00111001};
				  10'd110: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110000};
				  10'd111: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110001};
				  10'd112: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110010};
				  10'd113: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110011};
				  10'd114: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110100};
				  10'd115: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110101};
				  10'd116: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110110};
				  10'd117: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00110111};
				  10'd118: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00111000};
				  10'd119: reg_data_out_q <= {8'b00110001,8'b00110001,8'b00111001};
				  10'd120: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110000};
				  10'd121: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110001};
				  10'd122: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110010};
				  10'd123: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110011};
				  10'd124: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110100};
				  10'd125: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110101};
				  10'd125: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110101};
				  10'd126: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110110};
				  10'd127: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00110111};
				  10'd128: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00111000};
				  10'd129: reg_data_out_q <= {8'b00110001,8'b00110010,8'b00111001};
				  10'd130: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110000};
				  10'd131: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110001};
				  10'd132: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110010};
				  10'd133: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110011};
				  10'd134: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110100};
				  10'd135: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110101};
				  10'd136: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110110};
				  10'd137: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00110111};
				  10'd138: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00111000};
				  10'd139: reg_data_out_q <= {8'b00110001,8'b00110011,8'b00111001};
				  10'd140: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110000};
				  10'd141: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110001};
				  10'd142: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110010};
				  10'd143: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110011};
				  10'd144: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110100};
				  10'd145: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110101};
				  10'd146: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110110};
				  10'd147: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00110111};
				  10'd148: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00111000};
				  10'd149: reg_data_out_q <= {8'b00110001,8'b00110100,8'b00111001};
				  10'd150: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110000};
				  10'd151: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110001};
				  10'd152: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110010};
				  10'd153: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110011};
				  10'd154: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110100};
				  10'd155: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110101};
				  10'd156: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110110};
				  10'd157: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00110111};
				  10'd158: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00111000};
				  10'd159: reg_data_out_q <= {8'b00110001,8'b00110101,8'b00111001};
				  10'd160: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110000};
				  10'd161: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110001};
				  10'd162: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110010};
				  10'd163: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110011};
				  10'd164: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110100};
				  10'd165: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110101};
				  10'd166: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110110};
				  10'd166: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110110};
				  10'd167: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00110111};
				  10'd168: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00111000};
				  10'd169: reg_data_out_q <= {8'b00110001,8'b00110110,8'b00111001};
				  10'd170: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110000};
				  10'd171: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110001};
				  10'd172: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110010};
				  10'd173: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110011};
				  10'd174: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110100};
				  10'd175: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110101};
				  10'd176: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110110};
				  10'd177: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00110111};
				  10'd178: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00111000};
				  10'd179: reg_data_out_q <= {8'b00110001,8'b00110111,8'b00111001};
				  10'd180: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110000};
				  10'd181: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110001};
				  10'd182: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110010};
				  10'd183: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110011};
				  10'd184: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110100};
				  10'd185: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110101};
				  10'd186: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110110};
				  10'd187: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00110111};
				  10'd188: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00111000};
				  10'd189: reg_data_out_q <= {8'b00110001,8'b00111000,8'b00111001};
				  10'd190: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110000};
				  10'd191: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110001};
				  10'd192: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110010};
				  10'd193: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110011};
				  10'd194: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110100};
				  10'd195: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110101};
				  10'd196: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110110};
				  10'd197: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00110111};
				  10'd198: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00111000};
				  10'd199: reg_data_out_q <= {8'b00110001,8'b00111001,8'b00111001};
				  10'd200: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110000};
				  10'd201: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110001};
				  10'd202: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110010};
				  10'd203: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110011};
				  10'd204: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110100};
				  10'd205: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110101};
				  10'd206: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110110};
				  10'd207: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00110111};
				  10'd208: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00111000};
				  10'd208: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00111000};
				  10'd209: reg_data_out_q <= {8'b00110010,8'b00110000,8'b00111001};
				  10'd210: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110000};
				  10'd211: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110001};
				  10'd212: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110010};
				  10'd213: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110011};
				  10'd214: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110100};
				  10'd215: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110101};
				  10'd216: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110110};
				  10'd217: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00110111};
				  10'd218: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00111000};
				  10'd219: reg_data_out_q <= {8'b00110010,8'b00110001,8'b00111001};
				  10'd220: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110000};
				  10'd221: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110001};
				  10'd222: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110010};
				  10'd223: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110011};
				  10'd224: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110100};
				  10'd225: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110101};
				  10'd226: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110110};
				  10'd227: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00110111};
				  10'd228: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00111000};
				  10'd229: reg_data_out_q <= {8'b00110010,8'b00110010,8'b00111001};
				  10'd230: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110000};
				  10'd231: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110001};
				  10'd232: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110010};
				  10'd233: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110011};
				  10'd234: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110100};
				  10'd235: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110101};
				  10'd236: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110110};
				  10'd237: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00110111};
				  10'd238: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00111000};
				  10'd239: reg_data_out_q <= {8'b00110010,8'b00110011,8'b00111001};
				  10'd240: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110000};
				  10'd241: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110001};
				  10'd242: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110010};
				  10'd243: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110011};
				  10'd244: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110100};
				  10'd245: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110101};
				  10'd246: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110110};
				  10'd247: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00110111};
				  10'd248: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00111000};
				  10'd249: reg_data_out_q <= {8'b00110010,8'b00110100,8'b00111001};
				  10'd250: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00000000};
				  10'd250: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110000};
				  10'd251: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110001};
				  10'd252: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110010};
				  10'd253: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110011};
				  10'd254: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110100};
				  10'd255: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110101};
				  10'd256: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110110};
				  10'd257: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00110111};
				  10'd258: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00111000};
				  10'd259: reg_data_out_q <= {8'b00110010,8'b00110101,8'b00111001};
				  10'd260: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110000};
				  10'd261: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110001};
				  10'd262: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110010};
				  10'd263: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110011};
				  10'd264: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110100};
				  10'd265: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110101};
				  10'd266: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110110};
				  10'd267: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00110111};
				  10'd268: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00111000};
				  10'd269: reg_data_out_q <= {8'b00110010,8'b00110110,8'b00111001};
				  10'd270: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110000};
				  10'd271: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110001};
				  10'd272: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110010};
				  10'd273: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110011};
				  10'd274: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110100};
				  10'd275: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110101};
				  10'd276: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110110};
				  10'd277: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00110111};
				  10'd278: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00111000};
				  10'd279: reg_data_out_q <= {8'b00110010,8'b00110111,8'b00111001};
				  10'd280: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110000};
				  10'd281: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110001};
				  10'd282: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110010};
				  10'd283: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110011};
				  10'd284: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110100};
				  10'd285: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110101};
				  10'd286: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110110};
				  10'd287: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00110111};
				  10'd288: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00111000};
				  10'd289: reg_data_out_q <= {8'b00110010,8'b00111000,8'b00111001};
				  10'd290: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110000};
				  10'd291: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110001};
				  10'd291: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110001};
				  10'd292: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110010};
				  10'd293: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110011};
				  10'd294: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110100};
				  10'd295: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110101};
				  10'd296: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110110};
				  10'd297: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00110111};
				  10'd298: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00111000};
				  10'd299: reg_data_out_q <= {8'b00110010,8'b00111001,8'b00111001};
				  10'd300: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110000};
				  10'd301: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110001};
				  10'd302: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110010};
				  10'd303: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110011};
				  10'd304: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110100};
				  10'd305: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110101};
				  10'd306: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110110};
				  10'd307: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00110111};
				  10'd308: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00111000};
				  10'd309: reg_data_out_q <= {8'b00110011,8'b00110000,8'b00111001};
				  10'd310: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110000};
				  10'd311: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110001};
				  10'd312: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110010};
				  10'd313: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110011};
				  10'd314: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110100};
				  10'd315: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110101};
				  10'd316: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110110};
				  10'd317: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00110111};
				  10'd318: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00111000};
				  10'd319: reg_data_out_q <= {8'b00110011,8'b00110001,8'b00111001};
				  10'd320: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110000};
				  10'd321: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110001};
				  10'd322: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110010};
				  10'd323: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110011};
				  10'd324: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110100};
				  10'd325: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110101};
				  10'd326: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110110};
				  10'd327: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00110111};
				  10'd328: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00111000};
				  10'd329: reg_data_out_q <= {8'b00110011,8'b00110010,8'b00111001};
				  10'd330: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110000};
				  10'd331: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110001};
				  10'd332: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110010};
				  10'd333: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110011};
				  10'd333: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110011};
				  10'd334: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110100};
				  10'd335: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110101};
				  10'd336: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110110};
				  10'd337: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00110111};
				  10'd338: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00111000};
				  10'd339: reg_data_out_q <= {8'b00110011,8'b00110011,8'b00111001};
				  10'd340: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110000};
				  10'd341: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110001};
				  10'd342: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110010};
				  10'd343: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110011};
				  10'd344: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110100};
				  10'd345: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110101};
				  10'd346: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110110};
				  10'd347: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00110111};
				  10'd348: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00111000};
				  10'd349: reg_data_out_q <= {8'b00110011,8'b00110100,8'b00111001};
				  10'd350: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110000};
				  10'd351: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110001};
				  10'd352: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110010};
				  10'd353: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110011};
				  10'd354: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110100};
				  10'd355: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110101};
				  10'd356: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110110};
				  10'd357: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00110111};
				  10'd358: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00111000};
				  10'd359: reg_data_out_q <= {8'b00110011,8'b00110101,8'b00111001};
				  10'd360: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110000};
				  10'd361: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110001};
				  10'd362: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110010};
				  10'd363: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110011};
				  10'd364: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110100};
				  10'd365: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110101};
				  10'd366: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110110};
				  10'd367: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00110111};
				  10'd368: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00111000};
				  10'd369: reg_data_out_q <= {8'b00110011,8'b00110110,8'b00111001};
				  10'd370: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110000};
				  10'd371: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110001};
				  10'd372: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110010};
				  10'd373: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110011};
				  10'd374: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110100};
				  10'd375: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110101};
				  10'd375: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110101};
				  10'd376: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110110};
				  10'd377: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00110111};
				  10'd378: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00111000};
				  10'd379: reg_data_out_q <= {8'b00110011,8'b00110111,8'b00111001};
				  10'd380: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110000};
				  10'd381: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110001};
				  10'd382: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110010};
				  10'd383: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110011};
				  10'd384: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110100};
				  10'd385: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110101};
				  10'd386: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110110};
				  10'd387: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00110111};
				  10'd388: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00111000};
				  10'd389: reg_data_out_q <= {8'b00110011,8'b00111000,8'b00111001};
				  10'd390: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110000};
				  10'd391: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110001};
				  10'd392: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110010};
				  10'd393: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110011};
				  10'd394: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110100};
				  10'd395: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110101};
				  10'd396: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110110};
				  10'd397: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00110111};
				  10'd398: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00111000};
				  10'd399: reg_data_out_q <= {8'b00110011,8'b00111001,8'b00111001};
				  10'd400: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110000};
				  10'd401: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110001};
				  10'd402: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110010};
				  10'd403: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110011};
				  10'd404: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110100};
				  10'd405: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110101};
				  10'd406: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110110};
				  10'd407: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00110111};
				  10'd408: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00111000};
				  10'd409: reg_data_out_q <= {8'b00110100,8'b00110000,8'b00111001};
				  10'd410: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110000};
				  10'd411: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110001};
				  10'd412: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110010};
				  10'd413: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110011};
				  10'd414: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110100};
				  10'd415: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110101};
				  10'd416: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110110};
				  10'd416: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110110};
				  10'd417: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00110111};
				  10'd418: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00111000};
				  10'd419: reg_data_out_q <= {8'b00110100,8'b00110001,8'b00111001};
				  10'd420: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110000};
				  10'd421: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110001};
				  10'd422: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110010};
				  10'd423: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110011};
				  10'd424: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110100};
				  10'd425: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110101};
				  10'd426: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110110};
				  10'd427: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00110111};
				  10'd428: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00111000};
				  10'd429: reg_data_out_q <= {8'b00110100,8'b00110010,8'b00111001};
				  10'd430: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110000};
				  10'd431: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110001};
				  10'd432: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110010};
				  10'd433: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110011};
				  10'd434: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110100};
				  10'd435: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110101};
				  10'd436: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110110};
				  10'd437: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00110111};
				  10'd438: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00111000};
				  10'd439: reg_data_out_q <= {8'b00110100,8'b00110011,8'b00111001};
				  10'd440: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110000};
				  10'd441: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110001};
				  10'd442: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110010};
				  10'd443: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110011};
				  10'd444: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110100};
				  10'd445: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110101};
				  10'd446: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110110};
				  10'd447: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00110111};
				  10'd448: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00111000};
				  10'd449: reg_data_out_q <= {8'b00110100,8'b00110100,8'b00111001};
				  10'd450: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110000};
				  10'd451: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110001};
				  10'd452: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110010};
				  10'd453: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110011};
				  10'd454: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110100};
				  10'd455: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110101};
				  10'd456: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110110};
				  10'd457: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00110111};
				  10'd458: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00111000};
				  10'd458: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00111000};
				  10'd459: reg_data_out_q <= {8'b00110100,8'b00110101,8'b00111001};
				  10'd460: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110000};
				  10'd461: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110001};
				  10'd462: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110010};
				  10'd463: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110011};
				  10'd464: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110100};
				  10'd465: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110101};
				  10'd466: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110110};
				  10'd467: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00110111};
				  10'd468: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00111000};
				  10'd469: reg_data_out_q <= {8'b00110100,8'b00110110,8'b00111001};
				  10'd470: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110000};
				  10'd471: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110001};
				  10'd472: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110010};
				  10'd473: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110011};
				  10'd474: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110100};
				  10'd475: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110101};
				  10'd476: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110110};
				  10'd477: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00110111};
				  10'd478: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00111000};
				  10'd479: reg_data_out_q <= {8'b00110100,8'b00110111,8'b00111001};
				  10'd480: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110000};
				  10'd481: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110001};
				  10'd482: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110010};
				  10'd483: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110011};
				  10'd484: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110100};
				  10'd485: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110101};
				  10'd486: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110110};
				  10'd487: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00110111};
				  10'd488: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00111000};
				  10'd489: reg_data_out_q <= {8'b00110100,8'b00111000,8'b00111001};
				  10'd490: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110000};
				  10'd491: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110001};
				  10'd492: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110010};
				  10'd493: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110011};
				  10'd494: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110100};
				  10'd495: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110101};
				  10'd496: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110110};
				  10'd497: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00110111};
				  10'd498: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00111000};
				  10'd499: reg_data_out_q <= {8'b00110100,8'b00111001,8'b00111001};
				  10'd500: reg_data_out_q <= {8'b00110101,8'b00000000,8'b00000000};
				  10'd500: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110000};
				  10'd501: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110001};
				  10'd502: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110010};
				  10'd503: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110011};
				  10'd504: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110100};
				  10'd505: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110101};
				  10'd506: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110110};
				  10'd507: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00110111};
				  10'd508: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00111000};
				  10'd509: reg_data_out_q <= {8'b00110101,8'b00110000,8'b00111001};
				  10'd510: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110000};
				  10'd511: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110001};
				  10'd512: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110010};
				  10'd513: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110011};
				  10'd514: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110100};
				  10'd515: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110101};
				  10'd516: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110110};
				  10'd517: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00110111};
				  10'd518: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00111000};
				  10'd519: reg_data_out_q <= {8'b00110101,8'b00110001,8'b00111001};
				  10'd520: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110000};
				  10'd521: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110001};
				  10'd522: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110010};
				  10'd523: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110011};
				  10'd524: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110100};
				  10'd525: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110101};
				  10'd526: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110110};
				  10'd527: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00110111};
				  10'd528: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00111000};
				  10'd529: reg_data_out_q <= {8'b00110101,8'b00110010,8'b00111001};
				  10'd530: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110000};
				  10'd531: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110001};
				  10'd532: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110010};
				  10'd533: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110011};
				  10'd534: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110100};
				  10'd535: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110101};
				  10'd536: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110110};
				  10'd537: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00110111};
				  10'd538: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00111000};
				  10'd539: reg_data_out_q <= {8'b00110101,8'b00110011,8'b00111001};
				  10'd540: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110000};
				  10'd541: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110001};
				  10'd541: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110001};
				  10'd542: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110010};
				  10'd543: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110011};
				  10'd544: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110100};
				  10'd545: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110101};
				  10'd546: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110110};
				  10'd547: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00110111};
				  10'd548: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00111000};
				  10'd549: reg_data_out_q <= {8'b00110101,8'b00110100,8'b00111001};
				  10'd550: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110000};
				  10'd551: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110001};
				  10'd552: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110010};
				  10'd553: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110011};
				  10'd554: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110100};
				  10'd555: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110101};
				  10'd556: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110110};
				  10'd557: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00110111};
				  10'd558: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00111000};
				  10'd559: reg_data_out_q <= {8'b00110101,8'b00110101,8'b00111001};
				  10'd560: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110000};
				  10'd561: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110001};
				  10'd562: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110010};
				  10'd563: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110011};
				  10'd564: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110100};
				  10'd565: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110101};
				  10'd566: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110110};
				  10'd567: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00110111};
				  10'd568: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00111000};
				  10'd569: reg_data_out_q <= {8'b00110101,8'b00110110,8'b00111001};
				  10'd570: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110000};
				  10'd571: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110001};
				  10'd572: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110010};
				  10'd573: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110011};
				  10'd574: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110100};
				  10'd575: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110101};
				  10'd576: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110110};
				  10'd577: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00110111};
				  10'd578: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00111000};
				  10'd579: reg_data_out_q <= {8'b00110101,8'b00110111,8'b00111001};
				  10'd580: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110000};
				  10'd581: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110001};
				  10'd582: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110010};
				  10'd583: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110011};
				  10'd583: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110011};
				  10'd584: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110100};
				  10'd585: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110101};
				  10'd586: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110110};
				  10'd587: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00110111};
				  10'd588: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00111000};
				  10'd589: reg_data_out_q <= {8'b00110101,8'b00111000,8'b00111001};
				  10'd590: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110000};
				  10'd591: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110001};
				  10'd592: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110010};
				  10'd593: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110011};
				  10'd594: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110100};
				  10'd595: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110101};
				  10'd596: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110110};
				  10'd597: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00110111};
				  10'd598: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00111000};
				  10'd599: reg_data_out_q <= {8'b00110101,8'b00111001,8'b00111001};
				  10'd600: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110000};
				  10'd601: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110001};
				  10'd602: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110010};
				  10'd603: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110011};
				  10'd604: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110100};
				  10'd605: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110101};
				  10'd606: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110110};
				  10'd607: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00110111};
				  10'd608: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00111000};
				  10'd609: reg_data_out_q <= {8'b00110110,8'b00110000,8'b00111001};
				  10'd610: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110000};
				  10'd611: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110001};
				  10'd612: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110010};
				  10'd613: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110011};
				  10'd614: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110100};
				  10'd615: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110101};
				  10'd616: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110110};
				  10'd617: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00110111};
				  10'd618: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00111000};
				  10'd619: reg_data_out_q <= {8'b00110110,8'b00110001,8'b00111001};
				  10'd620: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110000};
				  10'd621: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110001};
				  10'd622: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110010};
				  10'd623: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110011};
				  10'd624: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110100};
				  10'd625: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110101};
				  10'd625: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110101};
				  10'd626: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110110};
				  10'd627: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00110111};
				  10'd628: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00111000};
				  10'd629: reg_data_out_q <= {8'b00110110,8'b00110010,8'b00111001};
				  10'd630: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110000};
				  10'd631: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110001};
				  10'd632: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110010};
				  10'd633: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110011};
				  10'd634: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110100};
				  10'd635: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110101};
				  10'd636: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110110};
				  10'd637: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00110111};
				  10'd638: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00111000};
				  10'd639: reg_data_out_q <= {8'b00110110,8'b00110011,8'b00111001};
				  10'd640: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110000};
				  10'd641: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110001};
				  10'd642: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110010};
				  10'd643: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110011};
				  10'd644: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110100};
				  10'd645: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110101};
				  10'd646: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110110};
				  10'd647: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00110111};
				  10'd648: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00111000};
				  10'd649: reg_data_out_q <= {8'b00110110,8'b00110100,8'b00111001};
				  10'd650: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110000};
				  10'd651: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110001};
				  10'd652: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110010};
				  10'd653: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110011};
				  10'd654: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110100};
				  10'd655: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110101};
				  10'd656: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110110};
				  10'd657: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00110111};
				  10'd658: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00111000};
				  10'd659: reg_data_out_q <= {8'b00110110,8'b00110101,8'b00111001};
				  10'd660: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110000};
				  10'd661: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110001};
				  10'd662: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110010};
				  10'd663: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110011};
				  10'd664: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110100};
				  10'd665: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110101};
				  10'd666: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110110};
				  10'd666: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110110};
				  10'd667: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00110111};
				  10'd668: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00111000};
				  10'd669: reg_data_out_q <= {8'b00110110,8'b00110110,8'b00111001};
				  10'd670: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110000};
				  10'd671: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110001};
				  10'd672: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110010};
				  10'd673: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110011};
				  10'd674: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110100};
				  10'd675: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110101};
				  10'd676: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110110};
				  10'd677: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00110111};
				  10'd678: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00111000};
				  10'd679: reg_data_out_q <= {8'b00110110,8'b00110111,8'b00111001};
				  10'd680: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110000};
				  10'd681: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110001};
				  10'd682: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110010};
				  10'd683: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110011};
				  10'd684: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110100};
				  10'd685: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110101};
				  10'd686: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110110};
				  10'd687: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00110111};
				  10'd688: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00111000};
				  10'd689: reg_data_out_q <= {8'b00110110,8'b00111000,8'b00111001};
				  10'd690: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110000};
				  10'd691: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110001};
				  10'd692: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110010};
				  10'd693: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110011};
				  10'd694: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110100};
				  10'd695: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110101};
				  10'd696: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110110};
				  10'd697: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00110111};
				  10'd698: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00111000};
				  10'd699: reg_data_out_q <= {8'b00110110,8'b00111001,8'b00111001};
				  10'd700: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110000};
				  10'd701: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110001};
				  10'd702: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110010};
				  10'd703: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110011};
				  10'd704: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110100};
				  10'd705: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110101};
				  10'd706: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110110};
				  10'd707: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00110111};
				  10'd708: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00111000};
				  10'd708: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00111000};
				  10'd709: reg_data_out_q <= {8'b00110111,8'b00110000,8'b00111001};
				  10'd710: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110000};
				  10'd711: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110001};
				  10'd712: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110010};
				  10'd713: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110011};
				  10'd714: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110100};
				  10'd715: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110101};
				  10'd716: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110110};
				  10'd717: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00110111};
				  10'd718: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00111000};
				  10'd719: reg_data_out_q <= {8'b00110111,8'b00110001,8'b00111001};
				  10'd720: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110000};
				  10'd721: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110001};
				  10'd722: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110010};
				  10'd723: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110011};
				  10'd724: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110100};
				  10'd725: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110101};
				  10'd726: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110110};
				  10'd727: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00110111};
				  10'd728: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00111000};
				  10'd729: reg_data_out_q <= {8'b00110111,8'b00110010,8'b00111001};
				  10'd730: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110000};
				  10'd731: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110001};
				  10'd732: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110010};
				  10'd733: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110011};
				  10'd734: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110100};
				  10'd735: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110101};
				  10'd736: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110110};
				  10'd737: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00110111};
				  10'd738: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00111000};
				  10'd739: reg_data_out_q <= {8'b00110111,8'b00110011,8'b00111001};
				  10'd740: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110000};
				  10'd741: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110001};
				  10'd742: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110010};
				  10'd743: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110011};
				  10'd744: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110100};
				  10'd745: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110101};
				  10'd746: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110110};
				  10'd747: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00110111};
				  10'd748: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00111000};
				  10'd749: reg_data_out_q <= {8'b00110111,8'b00110100,8'b00111001};
				  10'd750: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00000000};
				  10'd750: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110000};
				  10'd751: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110001};
				  10'd752: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110010};
				  10'd753: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110011};
				  10'd754: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110100};
				  10'd755: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110101};
				  10'd756: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110110};
				  10'd757: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00110111};
				  10'd758: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00111000};
				  10'd759: reg_data_out_q <= {8'b00110111,8'b00110101,8'b00111001};
				  10'd760: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110000};
				  10'd761: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110001};
				  10'd762: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110010};
				  10'd763: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110011};
				  10'd764: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110100};
				  10'd765: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110101};
				  10'd766: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110110};
				  10'd767: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00110111};
				  10'd768: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00111000};
				  10'd769: reg_data_out_q <= {8'b00110111,8'b00110110,8'b00111001};
				  10'd770: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110000};
				  10'd771: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110001};
				  10'd772: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110010};
				  10'd773: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110011};
				  10'd774: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110100};
				  10'd775: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110101};
				  10'd776: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110110};
				  10'd777: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00110111};
				  10'd778: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00111000};
				  10'd779: reg_data_out_q <= {8'b00110111,8'b00110111,8'b00111001};
				  10'd780: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110000};
				  10'd781: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110001};
				  10'd782: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110010};
				  10'd783: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110011};
				  10'd784: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110100};
				  10'd785: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110101};
				  10'd786: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110110};
				  10'd787: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00110111};
				  10'd788: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00111000};
				  10'd789: reg_data_out_q <= {8'b00110111,8'b00111000,8'b00111001};
				  10'd790: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110000};
				  10'd791: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110001};
				  10'd791: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110001};
				  10'd792: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110010};
				  10'd793: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110011};
				  10'd794: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110100};
				  10'd795: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110101};
				  10'd796: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110110};
				  10'd797: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00110111};
				  10'd798: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00111000};
				  10'd799: reg_data_out_q <= {8'b00110111,8'b00111001,8'b00111001};
				  10'd800: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110000};
				  10'd801: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110001};
				  10'd802: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110010};
				  10'd803: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110011};
				  10'd804: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110100};
				  10'd805: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110101};
				  10'd806: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110110};
				  10'd807: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00110111};
				  10'd808: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00111000};
				  10'd809: reg_data_out_q <= {8'b00111000,8'b00110000,8'b00111001};
				  10'd810: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110000};
				  10'd811: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110001};
				  10'd812: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110010};
				  10'd813: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110011};
				  10'd814: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110100};
				  10'd815: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110101};
				  10'd816: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110110};
				  10'd817: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00110111};
				  10'd818: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00111000};
				  10'd819: reg_data_out_q <= {8'b00111000,8'b00110001,8'b00111001};
				  10'd820: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110000};
				  10'd821: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110001};
				  10'd822: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110010};
				  10'd823: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110011};
				  10'd824: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110100};
				  10'd825: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110101};
				  10'd826: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110110};
				  10'd827: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00110111};
				  10'd828: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00111000};
				  10'd829: reg_data_out_q <= {8'b00111000,8'b00110010,8'b00111001};
				  10'd830: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110000};
				  10'd831: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110001};
				  10'd832: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110010};
				  10'd833: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110011};
				  10'd833: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110011};
				  10'd834: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110100};
				  10'd835: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110101};
				  10'd836: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110110};
				  10'd837: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00110111};
				  10'd838: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00111000};
				  10'd839: reg_data_out_q <= {8'b00111000,8'b00110011,8'b00111001};
				  10'd840: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110000};
				  10'd841: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110001};
				  10'd842: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110010};
				  10'd843: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110011};
				  10'd844: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110100};
				  10'd845: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110101};
				  10'd846: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110110};
				  10'd847: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00110111};
				  10'd848: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00111000};
				  10'd849: reg_data_out_q <= {8'b00111000,8'b00110100,8'b00111001};
				  10'd850: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110000};
				  10'd851: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110001};
				  10'd852: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110010};
				  10'd853: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110011};
				  10'd854: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110100};
				  10'd855: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110101};
				  10'd856: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110110};
				  10'd857: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00110111};
				  10'd858: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00111000};
				  10'd859: reg_data_out_q <= {8'b00111000,8'b00110101,8'b00111001};
				  10'd860: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110000};
				  10'd861: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110001};
				  10'd862: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110010};
				  10'd863: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110011};
				  10'd864: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110100};
				  10'd865: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110101};
				  10'd866: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110110};
				  10'd867: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00110111};
				  10'd868: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00111000};
				  10'd869: reg_data_out_q <= {8'b00111000,8'b00110110,8'b00111001};
				  10'd870: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110000};
				  10'd871: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110001};
				  10'd872: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110010};
				  10'd873: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110011};
				  10'd874: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110100};
				  10'd875: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110101};
				  10'd875: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110101};
				  10'd876: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110110};
				  10'd877: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00110111};
				  10'd878: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00111000};
				  10'd879: reg_data_out_q <= {8'b00111000,8'b00110111,8'b00111001};
				  10'd880: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110000};
				  10'd881: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110001};
				  10'd882: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110010};
				  10'd883: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110011};
				  10'd884: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110100};
				  10'd885: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110101};
				  10'd886: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110110};
				  10'd887: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00110111};
				  10'd888: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00111000};
				  10'd889: reg_data_out_q <= {8'b00111000,8'b00111000,8'b00111001};
				  10'd890: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110000};
				  10'd891: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110001};
				  10'd892: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110010};
				  10'd893: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110011};
				  10'd894: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110100};
				  10'd895: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110101};
				  10'd896: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110110};
				  10'd897: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00110111};
				  10'd898: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00111000};
				  10'd899: reg_data_out_q <= {8'b00111000,8'b00111001,8'b00111001};
				  10'd900: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110000};
				  10'd901: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110001};
				  10'd902: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110010};
				  10'd903: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110011};
				  10'd904: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110100};
				  10'd905: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110101};
				  10'd906: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110110};
				  10'd907: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00110111};
				  10'd908: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00111000};
				  10'd909: reg_data_out_q <= {8'b00111001,8'b00110000,8'b00111001};
				  10'd910: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110000};
				  10'd911: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110001};
				  10'd912: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110010};
				  10'd913: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110011};
				  10'd914: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110100};
				  10'd915: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110101};
				  10'd916: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110110};
				  10'd916: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110110};
				  10'd917: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00110111};
				  10'd918: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00111000};
				  10'd919: reg_data_out_q <= {8'b00111001,8'b00110001,8'b00111001};
				  10'd920: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110000};
				  10'd921: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110001};
				  10'd922: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110010};
				  10'd923: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110011};
				  10'd924: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110100};
				  10'd925: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110101};
				  10'd926: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110110};
				  10'd927: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00110111};
				  10'd928: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00111000};
				  10'd929: reg_data_out_q <= {8'b00111001,8'b00110010,8'b00111001};
				  10'd930: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110000};
				  10'd931: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110001};
				  10'd932: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110010};
				  10'd933: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110011};
				  10'd934: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110100};
				  10'd935: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110101};
				  10'd936: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110110};
				  10'd937: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00110111};
				  10'd938: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00111000};
				  10'd939: reg_data_out_q <= {8'b00111001,8'b00110011,8'b00111001};
				  10'd940: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110000};
				  10'd941: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110001};
				  10'd942: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110010};
				  10'd943: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110011};
				  10'd944: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110100};
				  10'd945: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110101};
				  10'd946: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110110};
				  10'd947: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00110111};
				  10'd948: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00111000};
				  10'd949: reg_data_out_q <= {8'b00111001,8'b00110100,8'b00111001};
				  10'd950: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110000};
				  10'd951: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110001};
				  10'd952: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110010};
				  10'd953: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110011};
				  10'd954: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110100};
				  10'd955: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110101};
				  10'd956: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110110};
				  10'd957: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00110111};
				  10'd958: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00111000};
				  10'd958: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00111000};
				  10'd959: reg_data_out_q <= {8'b00111001,8'b00110101,8'b00111001};
				  10'd960: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110000};
				  10'd961: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110001};
				  10'd962: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110010};
				  10'd963: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110011};
				  10'd964: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110100};
				  10'd965: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110101};
				  10'd966: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110110};
				  10'd967: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00110111};
				  10'd968: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00111000};
				  10'd969: reg_data_out_q <= {8'b00111001,8'b00110110,8'b00111001};
				  10'd970: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110000};
				  10'd971: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110001};
				  10'd972: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110010};
				  10'd973: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110011};
				  10'd974: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110100};
				  10'd975: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110101};
				  10'd976: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110110};
				  10'd977: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00110111};
				  10'd978: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00111000};
				  10'd979: reg_data_out_q <= {8'b00111001,8'b00110111,8'b00111001};
				  10'd980: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110000};
				  10'd981: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110001};
				  10'd982: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110010};
				  10'd983: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110011};
				  10'd984: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110100};
				  10'd985: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110101};
				  10'd986: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110110};
				  10'd987: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00110111};
				  10'd988: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00111000};
				  10'd989: reg_data_out_q <= {8'b00111001,8'b00111000,8'b00111001};
				  10'd990: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110000};
				  10'd991: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110001};
				  10'd992: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110010};
				  10'd993: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110011};
				  10'd994: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110100};
				  10'd995: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110101};
				  10'd996: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110110};
				  10'd997: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00110111};
				  10'd998: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00111000};
				  10'd999: reg_data_out_q <= {8'b00111001,8'b00111001,8'b00111001};
				  endcase
		end else begin
			if(again) begin
				reg_d_out_i <= 0;
				reg_data_out_q <=0;
			end
			reg_en_crc <=1'b0;
		end
	end

endmodule

