`define L_0 32'h5A000000
`define L_1 32'h35214E63
`define L_2 32'h1C128E80
`define L_3 32'h0E400224
`define L_4 32'h0727154C
`define L_5 32'h03946F29
`define L_6 32'h01CA5435
`define L_7 32'h00E52D8D
`define L_8 32'h007296C6
`define L_9 32'h00394B63
`define L_10 32'h001CA5B1
`define L_11 32'h000E52D8
`define L_12 32'h0007296C
`define L_13 32'h000394B6
`define L_14 32'h0001CA5B
`define L_15 32'h0000E52D
`define L_16 32'h00007296
`define L_17 32'h0000394B
`define L_18 32'h00001CA5
`define L_19 32'h00000E52
`define L_20 32'h00000729
`define L_21 32'h00000394
`define L_22 32'h000001CA
`define L_23 32'h000000E5
`define L_24 32'h00000072
`define L_25 32'h00000039
`define L_26 32'h0000001c
`define L_27 32'h0000000e
`define L_28 32'h00000007
`define L_29 32'h00000003
`define L_30 32'h00000001
`define L_31 32'h00000000

module atang(clk,en,rst,x_in,y_in,z_out,en_conv
    );
	 input clk,rst,en;
	 input  signed [31:0] x_in;
	 input  signed [31:0] y_in;
	 output [16:0] z_out;
	 //output [8:0] z_out;
	 output en_conv;

	 reg  signed [32:0] x_reg = 33'b0 ;
	 reg  signed [32:0] y_reg = 33'b0 ;
	 reg  [31:0] z_reg = 32'b0 ;
	 reg [3:0] state = 4'b0 ;
	 reg [5:0] count = 6'b0;
	 //reg [8:0] reg_aprx_z = 9'b0;
	 reg reg_en_conv=1'b0;
	 reg [9:0] reg_q = 10'b0;
	
	 parameter idle = 4'b0;
	 parameter start = 4'b0001;
	 parameter vect_mode = 4'b0010;
	 parameter end_state = 4'b0011;
	 parameter end_aproximari = 4'b0100;
	 parameter end_final = 4'b0101;
	 parameter final = 4'b0110;
	 
	 assign en_conv = reg_en_conv;
	 
	always @(posedge clk) begin
		case (state)
				idle : begin
					x_reg[32:0] <= 33'b0;
					y_reg[32:0] <= 33'b0;
					z_reg[31:0] <= 32'b0;
					//reg_aprx_z <=9'b0;
					count <= 6'b0;
					if (rst) 
						state <= idle;
					else
						state <= (en) ? start : idle ;
				end
				start: begin
					if (rst) 
						state <= idle;
					else begin
					x_reg[32:0] <= x_in[31:0] ;
					y_reg[32:0] <= y_in[31:0] ;
					state <= vect_mode ;
					end
				end
				vect_mode: begin
					if ( count[5:0] > 6'b011111 ) begin
						state <= end_final ;
						count <= 6'b0;
					end else begin
						x_reg[32:0] <= x_reg[32:0] + (d_sign ? -y_sift : y_sift);
						y_reg[32:0] <= (d_sign ? x_sift : -x_sift) + y_reg[32:0];
						z_reg[31:0] <= z_reg + (d_sign ? -unghi : unghi);
						count <= count + 1'b1 ;
						state <= vect_mode ;
					end
				end
				end_final : begin
					case(z_reg[24:15])
					  10'b0000000000: reg_q <= 10'd000;
					  10'b0000000001: reg_q <= 10'd000;
					  10'b0000000010: reg_q <= 10'd001;
					  10'b0000000011: reg_q <= 10'd002;
					  10'b0000000100: reg_q <= 10'd003;
					  10'b0000000101: reg_q <= 10'd004;
					  10'b0000000110: reg_q <= 10'd005;
					  10'b0000000111: reg_q <= 10'd006;
					  10'b0000001000: reg_q <= 10'd007;
					  10'b0000001001: reg_q <= 10'd008;
					  10'b0000001010: reg_q <= 10'd009;
					  10'b0000001011: reg_q <= 10'd010;
					  10'b0000001100: reg_q <= 10'd011;
					  10'b0000001101: reg_q <= 10'd012;
					  10'b0000001110: reg_q <= 10'd013;
					  10'b0000001111: reg_q <= 10'd014;
					  10'b0000010000: reg_q <= 10'd015;
					  10'b0000010001: reg_q <= 10'd016;
					  10'b0000010010: reg_q <= 10'd017;
					  10'b0000010011: reg_q <= 10'd018;
					  10'b0000010100: reg_q <= 10'd019;
					  10'b0000010101: reg_q <= 10'd020;
					  10'b0000010110: reg_q <= 10'd021;
					  10'b0000010111: reg_q <= 10'd022;
					  10'b0000011000: reg_q <= 10'd023;
					  10'b0000011001: reg_q <= 10'd024;
					  10'b0000011010: reg_q <= 10'd025;
					  10'b0000011011: reg_q <= 10'd026;
					  10'b0000011100: reg_q <= 10'd027;
					  10'b0000011101: reg_q <= 10'd028;
					  10'b0000011110: reg_q <= 10'd029;
					  10'b0000011111: reg_q <= 10'd030;
					  10'b0000100000: reg_q <= 10'd031;
					  10'b0000100001: reg_q <= 10'd032;
					  10'b0000100010: reg_q <= 10'd033;
					  10'b0000100011: reg_q <= 10'd034;
					  10'b0000100100: reg_q <= 10'd035;
					  10'b0000100101: reg_q <= 10'd036;
					  10'b0000100110: reg_q <= 10'd037;
					  10'b0000100111: reg_q <= 10'd038;
					  10'b0000101000: reg_q <= 10'd039;
					  10'b0000101001: reg_q <= 10'd040;
					  10'b0000101010: reg_q <= 10'd041;
					  10'b0000101011: reg_q <= 10'd041;
					  10'b0000101100: reg_q <= 10'd042;
					  10'b0000101101: reg_q <= 10'd043;
					  10'b0000101110: reg_q <= 10'd044;
					  10'b0000101111: reg_q <= 10'd045;
					  10'b0000110000: reg_q <= 10'd046;
					  10'b0000110001: reg_q <= 10'd047;
					  10'b0000110010: reg_q <= 10'd048;
					  10'b0000110011: reg_q <= 10'd049;
					  10'b0000110100: reg_q <= 10'd050;
					  10'b0000110101: reg_q <= 10'd051;
					  10'b0000110110: reg_q <= 10'd052;
					  10'b0000110111: reg_q <= 10'd053;
					  10'b0000111000: reg_q <= 10'd054;
					  10'b0000111001: reg_q <= 10'd055;
					  10'b0000111010: reg_q <= 10'd056;
					  10'b0000111011: reg_q <= 10'd057;
					  10'b0000111100: reg_q <= 10'd058;
					  10'b0000111101: reg_q <= 10'd059;
					  10'b0000111110: reg_q <= 10'd060;
					  10'b0000111111: reg_q <= 10'd061;
					  10'b0001000000: reg_q <= 10'd062;
					  10'b0001000001: reg_q <= 10'd063;
					  10'b0001000010: reg_q <= 10'd064;
					  10'b0001000011: reg_q <= 10'd065;
					  10'b0001000100: reg_q <= 10'd066;
					  10'b0001000101: reg_q <= 10'd067;
					  10'b0001000110: reg_q <= 10'd068;
					  10'b0001000111: reg_q <= 10'd069;
					  10'b0001001000: reg_q <= 10'd070;
					  10'b0001001001: reg_q <= 10'd071;
					  10'b0001001010: reg_q <= 10'd072;
					  10'b0001001011: reg_q <= 10'd073;
					  10'b0001001100: reg_q <= 10'd074;
					  10'b0001001101: reg_q <= 10'd075;
					  10'b0001001110: reg_q <= 10'd076;
					  10'b0001001111: reg_q <= 10'd077;
					  10'b0001010000: reg_q <= 10'd078;
					  10'b0001010001: reg_q <= 10'd079;
					  10'b0001010010: reg_q <= 10'd080;
					  10'b0001010011: reg_q <= 10'd081;
					  10'b0001010100: reg_q <= 10'd082;
					  10'b0001010101: reg_q <= 10'd083;
					  10'b0001010110: reg_q <= 10'd083;
					  10'b0001010111: reg_q <= 10'd084;
					  10'b0001011000: reg_q <= 10'd085;
					  10'b0001011001: reg_q <= 10'd086;
					  10'b0001011010: reg_q <= 10'd087;
					  10'b0001011011: reg_q <= 10'd088;
					  10'b0001011100: reg_q <= 10'd089;
					  10'b0001011101: reg_q <= 10'd090;
					  10'b0001011110: reg_q <= 10'd091;
					  10'b0001011111: reg_q <= 10'd092;
					  10'b0001100000: reg_q <= 10'd093;
					  10'b0001100001: reg_q <= 10'd094;
					  10'b0001100010: reg_q <= 10'd095;
					  10'b0001100011: reg_q <= 10'd096;
					  10'b0001100100: reg_q <= 10'd097;
					  10'b0001100101: reg_q <= 10'd098;
					  10'b0001100110: reg_q <= 10'd099;
					  10'b0001100111: reg_q <= 10'd100;
					  10'b0001101000: reg_q <= 10'd101;
					  10'b0001101001: reg_q <= 10'd102;
					  10'b0001101010: reg_q <= 10'd103;
					  10'b0001101011: reg_q <= 10'd104;
					  10'b0001101100: reg_q <= 10'd105;
					  10'b0001101101: reg_q <= 10'd106;
					  10'b0001101110: reg_q <= 10'd107;
					  10'b0001101111: reg_q <= 10'd108;
					  10'b0001110000: reg_q <= 10'd109;
					  10'b0001110001: reg_q <= 10'd110;
					  10'b0001110010: reg_q <= 10'd111;
					  10'b0001110011: reg_q <= 10'd112;
					  10'b0001110100: reg_q <= 10'd113;
					  10'b0001110101: reg_q <= 10'd114;
					  10'b0001110110: reg_q <= 10'd115;
					  10'b0001110111: reg_q <= 10'd116;
					  10'b0001111000: reg_q <= 10'd117;
					  10'b0001111001: reg_q <= 10'd118;
					  10'b0001111010: reg_q <= 10'd119;
					  10'b0001111011: reg_q <= 10'd120;
					  10'b0001111100: reg_q <= 10'd121;
					  10'b0001111101: reg_q <= 10'd122;
					  10'b0001111110: reg_q <= 10'd123;
					  10'b0001111111: reg_q <= 10'd124;
					  10'b0010000000: reg_q <= 10'd125;
					  10'b0010000001: reg_q <= 10'd125;
					  10'b0010000010: reg_q <= 10'd126;
					  10'b0010000011: reg_q <= 10'd127;
					  10'b0010000100: reg_q <= 10'd128;
					  10'b0010000101: reg_q <= 10'd129;
					  10'b0010000110: reg_q <= 10'd130;
					  10'b0010000111: reg_q <= 10'd131;
					  10'b0010001000: reg_q <= 10'd132;
					  10'b0010001001: reg_q <= 10'd133;
					  10'b0010001010: reg_q <= 10'd134;
					  10'b0010001011: reg_q <= 10'd135;
					  10'b0010001100: reg_q <= 10'd136;
					  10'b0010001101: reg_q <= 10'd137;
					  10'b0010001110: reg_q <= 10'd138;
					  10'b0010001111: reg_q <= 10'd139;
					  10'b0010010000: reg_q <= 10'd140;
					  10'b0010010001: reg_q <= 10'd141;
					  10'b0010010010: reg_q <= 10'd142;
					  10'b0010010011: reg_q <= 10'd143;
					  10'b0010010100: reg_q <= 10'd144;
					  10'b0010010101: reg_q <= 10'd145;
					  10'b0010010110: reg_q <= 10'd146;
					  10'b0010010111: reg_q <= 10'd147;
					  10'b0010011000: reg_q <= 10'd148;
					  10'b0010011001: reg_q <= 10'd149;
					  10'b0010011010: reg_q <= 10'd150;
					  10'b0010011011: reg_q <= 10'd151;
					  10'b0010011100: reg_q <= 10'd152;
					  10'b0010011101: reg_q <= 10'd153;
					  10'b0010011110: reg_q <= 10'd154;
					  10'b0010011111: reg_q <= 10'd155;
					  10'b0010100000: reg_q <= 10'd156;
					  10'b0010100001: reg_q <= 10'd157;
					  10'b0010100010: reg_q <= 10'd158;
					  10'b0010100011: reg_q <= 10'd159;
					  10'b0010100100: reg_q <= 10'd160;
					  10'b0010100101: reg_q <= 10'd161;
					  10'b0010100110: reg_q <= 10'd162;
					  10'b0010100111: reg_q <= 10'd163;
					  10'b0010101000: reg_q <= 10'd164;
					  10'b0010101001: reg_q <= 10'd165;
					  10'b0010101010: reg_q <= 10'd166;
					  10'b0010101011: reg_q <= 10'd166;
					  10'b0010101100: reg_q <= 10'd167;
					  10'b0010101101: reg_q <= 10'd168;
					  10'b0010101110: reg_q <= 10'd169;
					  10'b0010101111: reg_q <= 10'd170;
					  10'b0010110000: reg_q <= 10'd171;
					  10'b0010110001: reg_q <= 10'd172;
					  10'b0010110010: reg_q <= 10'd173;
					  10'b0010110011: reg_q <= 10'd174;
					  10'b0010110100: reg_q <= 10'd175;
					  10'b0010110101: reg_q <= 10'd176;
					  10'b0010110110: reg_q <= 10'd177;
					  10'b0010110111: reg_q <= 10'd178;
					  10'b0010111000: reg_q <= 10'd179;
					  10'b0010111001: reg_q <= 10'd180;
					  10'b0010111010: reg_q <= 10'd181;
					  10'b0010111011: reg_q <= 10'd182;
					  10'b0010111100: reg_q <= 10'd183;
					  10'b0010111101: reg_q <= 10'd184;
					  10'b0010111110: reg_q <= 10'd185;
					  10'b0010111111: reg_q <= 10'd186;
					  10'b0011000000: reg_q <= 10'd187;
					  10'b0011000001: reg_q <= 10'd188;
					  10'b0011000010: reg_q <= 10'd189;
					  10'b0011000011: reg_q <= 10'd190;
					  10'b0011000100: reg_q <= 10'd191;
					  10'b0011000101: reg_q <= 10'd192;
					  10'b0011000110: reg_q <= 10'd193;
					  10'b0011000111: reg_q <= 10'd194;
					  10'b0011001000: reg_q <= 10'd195;
					  10'b0011001001: reg_q <= 10'd196;
					  10'b0011001010: reg_q <= 10'd197;
					  10'b0011001011: reg_q <= 10'd198;
					  10'b0011001100: reg_q <= 10'd199;
					  10'b0011001101: reg_q <= 10'd200;
					  10'b0011001110: reg_q <= 10'd201;
					  10'b0011001111: reg_q <= 10'd202;
					  10'b0011010000: reg_q <= 10'd203;
					  10'b0011010001: reg_q <= 10'd204;
					  10'b0011010010: reg_q <= 10'd205;
					  10'b0011010011: reg_q <= 10'd206;
					  10'b0011010100: reg_q <= 10'd207;
					  10'b0011010101: reg_q <= 10'd208;
					  10'b0011010110: reg_q <= 10'd208;
					  10'b0011010111: reg_q <= 10'd209;
					  10'b0011011000: reg_q <= 10'd210;
					  10'b0011011001: reg_q <= 10'd211;
					  10'b0011011010: reg_q <= 10'd212;
					  10'b0011011011: reg_q <= 10'd213;
					  10'b0011011100: reg_q <= 10'd214;
					  10'b0011011101: reg_q <= 10'd215;
					  10'b0011011110: reg_q <= 10'd216;
					  10'b0011011111: reg_q <= 10'd217;
					  10'b0011100000: reg_q <= 10'd218;
					  10'b0011100001: reg_q <= 10'd219;
					  10'b0011100010: reg_q <= 10'd220;
					  10'b0011100011: reg_q <= 10'd221;
					  10'b0011100100: reg_q <= 10'd222;
					  10'b0011100101: reg_q <= 10'd223;
					  10'b0011100110: reg_q <= 10'd224;
					  10'b0011100111: reg_q <= 10'd225;
					  10'b0011101000: reg_q <= 10'd226;
					  10'b0011101001: reg_q <= 10'd227;
					  10'b0011101010: reg_q <= 10'd228;
					  10'b0011101011: reg_q <= 10'd229;
					  10'b0011101100: reg_q <= 10'd230;
					  10'b0011101101: reg_q <= 10'd231;
					  10'b0011101110: reg_q <= 10'd232;
					  10'b0011101111: reg_q <= 10'd233;
					  10'b0011110000: reg_q <= 10'd234;
					  10'b0011110001: reg_q <= 10'd235;
					  10'b0011110010: reg_q <= 10'd236;
					  10'b0011110011: reg_q <= 10'd237;
					  10'b0011110100: reg_q <= 10'd238;
					  10'b0011110101: reg_q <= 10'd239;
					  10'b0011110110: reg_q <= 10'd240;
					  10'b0011110111: reg_q <= 10'd241;
					  10'b0011111000: reg_q <= 10'd242;
					  10'b0011111001: reg_q <= 10'd243;
					  10'b0011111010: reg_q <= 10'd244;
					  10'b0011111011: reg_q <= 10'd245;
					  10'b0011111100: reg_q <= 10'd246;
					  10'b0011111101: reg_q <= 10'd247;
					  10'b0011111110: reg_q <= 10'd248;
					  10'b0011111111: reg_q <= 10'd249;
					  10'b0100000000: reg_q <= 10'd250;
					  10'b0100000001: reg_q <= 10'd250;
					  10'b0100000010: reg_q <= 10'd251;
					  10'b0100000011: reg_q <= 10'd252;
					  10'b0100000100: reg_q <= 10'd253;
					  10'b0100000101: reg_q <= 10'd254;
					  10'b0100000110: reg_q <= 10'd255;
					  10'b0100000111: reg_q <= 10'd256;
					  10'b0100001000: reg_q <= 10'd257;
					  10'b0100001001: reg_q <= 10'd258;
					  10'b0100001010: reg_q <= 10'd259;
					  10'b0100001011: reg_q <= 10'd260;
					  10'b0100001100: reg_q <= 10'd261;
					  10'b0100001101: reg_q <= 10'd262;
					  10'b0100001110: reg_q <= 10'd263;
					  10'b0100001111: reg_q <= 10'd264;
					  10'b0100010000: reg_q <= 10'd265;
					  10'b0100010001: reg_q <= 10'd266;
					  10'b0100010010: reg_q <= 10'd267;
					  10'b0100010011: reg_q <= 10'd268;
					  10'b0100010100: reg_q <= 10'd269;
					  10'b0100010101: reg_q <= 10'd270;
					  10'b0100010110: reg_q <= 10'd271;
					  10'b0100010111: reg_q <= 10'd272;
					  10'b0100011000: reg_q <= 10'd273;
					  10'b0100011001: reg_q <= 10'd274;
					  10'b0100011010: reg_q <= 10'd275;
					  10'b0100011011: reg_q <= 10'd276;
					  10'b0100011100: reg_q <= 10'd277;
					  10'b0100011101: reg_q <= 10'd278;
					  10'b0100011110: reg_q <= 10'd279;
					  10'b0100011111: reg_q <= 10'd280;
					  10'b0100100000: reg_q <= 10'd281;
					  10'b0100100001: reg_q <= 10'd282;
					  10'b0100100010: reg_q <= 10'd283;
					  10'b0100100011: reg_q <= 10'd284;
					  10'b0100100100: reg_q <= 10'd285;
					  10'b0100100101: reg_q <= 10'd286;
					  10'b0100100110: reg_q <= 10'd287;
					  10'b0100100111: reg_q <= 10'd288;
					  10'b0100101000: reg_q <= 10'd289;
					  10'b0100101001: reg_q <= 10'd290;
					  10'b0100101010: reg_q <= 10'd291;
					  10'b0100101011: reg_q <= 10'd291;
					  10'b0100101100: reg_q <= 10'd292;
					  10'b0100101101: reg_q <= 10'd293;
					  10'b0100101110: reg_q <= 10'd294;
					  10'b0100101111: reg_q <= 10'd295;
					  10'b0100110000: reg_q <= 10'd296;
					  10'b0100110001: reg_q <= 10'd297;
					  10'b0100110010: reg_q <= 10'd298;
					  10'b0100110011: reg_q <= 10'd299;
					  10'b0100110100: reg_q <= 10'd300;
					  10'b0100110101: reg_q <= 10'd301;
					  10'b0100110110: reg_q <= 10'd302;
					  10'b0100110111: reg_q <= 10'd303;
					  10'b0100111000: reg_q <= 10'd304;
					  10'b0100111001: reg_q <= 10'd305;
					  10'b0100111010: reg_q <= 10'd306;
					  10'b0100111011: reg_q <= 10'd307;
					  10'b0100111100: reg_q <= 10'd308;
					  10'b0100111101: reg_q <= 10'd309;
					  10'b0100111110: reg_q <= 10'd310;
					  10'b0100111111: reg_q <= 10'd311;
					  10'b0101000000: reg_q <= 10'd312;
					  10'b0101000001: reg_q <= 10'd313;
					  10'b0101000010: reg_q <= 10'd314;
					  10'b0101000011: reg_q <= 10'd315;
					  10'b0101000100: reg_q <= 10'd316;
					  10'b0101000101: reg_q <= 10'd317;
					  10'b0101000110: reg_q <= 10'd318;
					  10'b0101000111: reg_q <= 10'd319;
					  10'b0101001000: reg_q <= 10'd320;
					  10'b0101001001: reg_q <= 10'd321;
					  10'b0101001010: reg_q <= 10'd322;
					  10'b0101001011: reg_q <= 10'd323;
					  10'b0101001100: reg_q <= 10'd324;
					  10'b0101001101: reg_q <= 10'd325;
					  10'b0101001110: reg_q <= 10'd326;
					  10'b0101001111: reg_q <= 10'd327;
					  10'b0101010000: reg_q <= 10'd328;
					  10'b0101010001: reg_q <= 10'd329;
					  10'b0101010010: reg_q <= 10'd330;
					  10'b0101010011: reg_q <= 10'd331;
					  10'b0101010100: reg_q <= 10'd332;
					  10'b0101010101: reg_q <= 10'd333;
					  10'b0101010110: reg_q <= 10'd333;
					  10'b0101010111: reg_q <= 10'd334;
					  10'b0101011000: reg_q <= 10'd335;
					  10'b0101011001: reg_q <= 10'd336;
					  10'b0101011010: reg_q <= 10'd337;
					  10'b0101011011: reg_q <= 10'd338;
					  10'b0101011100: reg_q <= 10'd339;
					  10'b0101011101: reg_q <= 10'd340;
					  10'b0101011110: reg_q <= 10'd341;
					  10'b0101011111: reg_q <= 10'd342;
					  10'b0101100000: reg_q <= 10'd343;
					  10'b0101100001: reg_q <= 10'd344;
					  10'b0101100010: reg_q <= 10'd345;
					  10'b0101100011: reg_q <= 10'd346;
					  10'b0101100100: reg_q <= 10'd347;
					  10'b0101100101: reg_q <= 10'd348;
					  10'b0101100110: reg_q <= 10'd349;
					  10'b0101100111: reg_q <= 10'd350;
					  10'b0101101000: reg_q <= 10'd351;
					  10'b0101101001: reg_q <= 10'd352;
					  10'b0101101010: reg_q <= 10'd353;
					  10'b0101101011: reg_q <= 10'd354;
					  10'b0101101100: reg_q <= 10'd355;
					  10'b0101101101: reg_q <= 10'd356;
					  10'b0101101110: reg_q <= 10'd357;
					  10'b0101101111: reg_q <= 10'd358;
					  10'b0101110000: reg_q <= 10'd359;
					  10'b0101110001: reg_q <= 10'd360;
					  10'b0101110010: reg_q <= 10'd361;
					  10'b0101110011: reg_q <= 10'd362;
					  10'b0101110100: reg_q <= 10'd363;
					  10'b0101110101: reg_q <= 10'd364;
					  10'b0101110110: reg_q <= 10'd365;
					  10'b0101110111: reg_q <= 10'd366;
					  10'b0101111000: reg_q <= 10'd367;
					  10'b0101111001: reg_q <= 10'd368;
					  10'b0101111010: reg_q <= 10'd369;
					  10'b0101111011: reg_q <= 10'd370;
					  10'b0101111100: reg_q <= 10'd371;
					  10'b0101111101: reg_q <= 10'd372;
					  10'b0101111110: reg_q <= 10'd373;
					  10'b0101111111: reg_q <= 10'd374;
					  10'b0110000000: reg_q <= 10'd375;
					  10'b0110000001: reg_q <= 10'd375;
					  10'b0110000010: reg_q <= 10'd376;
					  10'b0110000011: reg_q <= 10'd377;
					  10'b0110000100: reg_q <= 10'd378;
					  10'b0110000101: reg_q <= 10'd379;
					  10'b0110000110: reg_q <= 10'd380;
					  10'b0110000111: reg_q <= 10'd381;
					  10'b0110001000: reg_q <= 10'd382;
					  10'b0110001001: reg_q <= 10'd383;
					  10'b0110001010: reg_q <= 10'd384;
					  10'b0110001011: reg_q <= 10'd385;
					  10'b0110001100: reg_q <= 10'd386;
					  10'b0110001101: reg_q <= 10'd387;
					  10'b0110001110: reg_q <= 10'd388;
					  10'b0110001111: reg_q <= 10'd389;
					  10'b0110010000: reg_q <= 10'd390;
					  10'b0110010001: reg_q <= 10'd391;
					  10'b0110010010: reg_q <= 10'd392;
					  10'b0110010011: reg_q <= 10'd393;
					  10'b0110010100: reg_q <= 10'd394;
					  10'b0110010101: reg_q <= 10'd395;
					  10'b0110010110: reg_q <= 10'd396;
					  10'b0110010111: reg_q <= 10'd397;
					  10'b0110011000: reg_q <= 10'd398;
					  10'b0110011001: reg_q <= 10'd399;
					  10'b0110011010: reg_q <= 10'd400;
					  10'b0110011011: reg_q <= 10'd401;
					  10'b0110011100: reg_q <= 10'd402;
					  10'b0110011101: reg_q <= 10'd403;
					  10'b0110011110: reg_q <= 10'd404;
					  10'b0110011111: reg_q <= 10'd405;
					  10'b0110100000: reg_q <= 10'd406;
					  10'b0110100001: reg_q <= 10'd407;
					  10'b0110100010: reg_q <= 10'd408;
					  10'b0110100011: reg_q <= 10'd409;
					  10'b0110100100: reg_q <= 10'd410;
					  10'b0110100101: reg_q <= 10'd411;
					  10'b0110100110: reg_q <= 10'd412;
					  10'b0110100111: reg_q <= 10'd413;
					  10'b0110101000: reg_q <= 10'd414;
					  10'b0110101001: reg_q <= 10'd415;
					  10'b0110101010: reg_q <= 10'd416;
					  10'b0110101011: reg_q <= 10'd416;
					  10'b0110101100: reg_q <= 10'd417;
					  10'b0110101101: reg_q <= 10'd418;
					  10'b0110101110: reg_q <= 10'd419;
					  10'b0110101111: reg_q <= 10'd420;
					  10'b0110110000: reg_q <= 10'd421;
					  10'b0110110001: reg_q <= 10'd422;
					  10'b0110110010: reg_q <= 10'd423;
					  10'b0110110011: reg_q <= 10'd424;
					  10'b0110110100: reg_q <= 10'd425;
					  10'b0110110101: reg_q <= 10'd426;
					  10'b0110110110: reg_q <= 10'd427;
					  10'b0110110111: reg_q <= 10'd428;
					  10'b0110111000: reg_q <= 10'd429;
					  10'b0110111001: reg_q <= 10'd430;
					  10'b0110111010: reg_q <= 10'd431;
					  10'b0110111011: reg_q <= 10'd432;
					  10'b0110111100: reg_q <= 10'd433;
					  10'b0110111101: reg_q <= 10'd434;
					  10'b0110111110: reg_q <= 10'd435;
					  10'b0110111111: reg_q <= 10'd436;
					  10'b0111000000: reg_q <= 10'd437;
					  10'b0111000001: reg_q <= 10'd438;
					  10'b0111000010: reg_q <= 10'd439;
					  10'b0111000011: reg_q <= 10'd440;
					  10'b0111000100: reg_q <= 10'd441;
					  10'b0111000101: reg_q <= 10'd442;
					  10'b0111000110: reg_q <= 10'd443;
					  10'b0111000111: reg_q <= 10'd444;
					  10'b0111001000: reg_q <= 10'd445;
					  10'b0111001001: reg_q <= 10'd446;
					  10'b0111001010: reg_q <= 10'd447;
					  10'b0111001011: reg_q <= 10'd448;
					  10'b0111001100: reg_q <= 10'd449;
					  10'b0111001101: reg_q <= 10'd450;
					  10'b0111001110: reg_q <= 10'd451;
					  10'b0111001111: reg_q <= 10'd452;
					  10'b0111010000: reg_q <= 10'd453;
					  10'b0111010001: reg_q <= 10'd454;
					  10'b0111010010: reg_q <= 10'd455;
					  10'b0111010011: reg_q <= 10'd456;
					  10'b0111010100: reg_q <= 10'd457;
					  10'b0111010101: reg_q <= 10'd458;
					  10'b0111010110: reg_q <= 10'd458;
					  10'b0111010111: reg_q <= 10'd459;
					  10'b0111011000: reg_q <= 10'd460;
					  10'b0111011001: reg_q <= 10'd461;
					  10'b0111011010: reg_q <= 10'd462;
					  10'b0111011011: reg_q <= 10'd463;
					  10'b0111011100: reg_q <= 10'd464;
					  10'b0111011101: reg_q <= 10'd465;
					  10'b0111011110: reg_q <= 10'd466;
					  10'b0111011111: reg_q <= 10'd467;
					  10'b0111100000: reg_q <= 10'd468;
					  10'b0111100001: reg_q <= 10'd469;
					  10'b0111100010: reg_q <= 10'd470;
					  10'b0111100011: reg_q <= 10'd471;
					  10'b0111100100: reg_q <= 10'd472;
					  10'b0111100101: reg_q <= 10'd473;
					  10'b0111100110: reg_q <= 10'd474;
					  10'b0111100111: reg_q <= 10'd475;
					  10'b0111101000: reg_q <= 10'd476;
					  10'b0111101001: reg_q <= 10'd477;
					  10'b0111101010: reg_q <= 10'd478;
					  10'b0111101011: reg_q <= 10'd479;
					  10'b0111101100: reg_q <= 10'd480;
					  10'b0111101101: reg_q <= 10'd481;
					  10'b0111101110: reg_q <= 10'd482;
					  10'b0111101111: reg_q <= 10'd483;
					  10'b0111110000: reg_q <= 10'd484;
					  10'b0111110001: reg_q <= 10'd485;
					  10'b0111110010: reg_q <= 10'd486;
					  10'b0111110011: reg_q <= 10'd487;
					  10'b0111110100: reg_q <= 10'd488;
					  10'b0111110101: reg_q <= 10'd489;
					  10'b0111110110: reg_q <= 10'd490;
					  10'b0111110111: reg_q <= 10'd491;
					  10'b0111111000: reg_q <= 10'd492;
					  10'b0111111001: reg_q <= 10'd493;
					  10'b0111111010: reg_q <= 10'd494;
					  10'b0111111011: reg_q <= 10'd495;
					  10'b0111111100: reg_q <= 10'd496;
					  10'b0111111101: reg_q <= 10'd497;
					  10'b0111111110: reg_q <= 10'd498;
					  10'b0111111111: reg_q <= 10'd499;
					  10'b1000000000: reg_q <= 10'd500;
					  10'b1000000001: reg_q <= 10'd500;
					  10'b1000000010: reg_q <= 10'd501;
					  10'b1000000011: reg_q <= 10'd502;
					  10'b1000000100: reg_q <= 10'd503;
					  10'b1000000101: reg_q <= 10'd504;
					  10'b1000000110: reg_q <= 10'd505;
					  10'b1000000111: reg_q <= 10'd506;
					  10'b1000001000: reg_q <= 10'd507;
					  10'b1000001001: reg_q <= 10'd508;
					  10'b1000001010: reg_q <= 10'd509;
					  10'b1000001011: reg_q <= 10'd510;
					  10'b1000001100: reg_q <= 10'd511;
					  10'b1000001101: reg_q <= 10'd512;
					  10'b1000001110: reg_q <= 10'd513;
					  10'b1000001111: reg_q <= 10'd514;
					  10'b1000010000: reg_q <= 10'd515;
					  10'b1000010001: reg_q <= 10'd516;
					  10'b1000010010: reg_q <= 10'd517;
					  10'b1000010011: reg_q <= 10'd518;
					  10'b1000010100: reg_q <= 10'd519;
					  10'b1000010101: reg_q <= 10'd520;
					  10'b1000010110: reg_q <= 10'd521;
					  10'b1000010111: reg_q <= 10'd522;
					  10'b1000011000: reg_q <= 10'd523;
					  10'b1000011001: reg_q <= 10'd524;
					  10'b1000011010: reg_q <= 10'd525;
					  10'b1000011011: reg_q <= 10'd526;
					  10'b1000011100: reg_q <= 10'd527;
					  10'b1000011101: reg_q <= 10'd528;
					  10'b1000011110: reg_q <= 10'd529;
					  10'b1000011111: reg_q <= 10'd530;
					  10'b1000100000: reg_q <= 10'd531;
					  10'b1000100001: reg_q <= 10'd532;
					  10'b1000100010: reg_q <= 10'd533;
					  10'b1000100011: reg_q <= 10'd534;
					  10'b1000100100: reg_q <= 10'd535;
					  10'b1000100101: reg_q <= 10'd536;
					  10'b1000100110: reg_q <= 10'd537;
					  10'b1000100111: reg_q <= 10'd538;
					  10'b1000101000: reg_q <= 10'd539;
					  10'b1000101001: reg_q <= 10'd540;
					  10'b1000101010: reg_q <= 10'd541;
					  10'b1000101011: reg_q <= 10'd541;
					  10'b1000101100: reg_q <= 10'd542;
					  10'b1000101101: reg_q <= 10'd543;
					  10'b1000101110: reg_q <= 10'd544;
					  10'b1000101111: reg_q <= 10'd545;
					  10'b1000110000: reg_q <= 10'd546;
					  10'b1000110001: reg_q <= 10'd547;
					  10'b1000110010: reg_q <= 10'd548;
					  10'b1000110011: reg_q <= 10'd549;
					  10'b1000110100: reg_q <= 10'd550;
					  10'b1000110101: reg_q <= 10'd551;
					  10'b1000110110: reg_q <= 10'd552;
					  10'b1000110111: reg_q <= 10'd553;
					  10'b1000111000: reg_q <= 10'd554;
					  10'b1000111001: reg_q <= 10'd555;
					  10'b1000111010: reg_q <= 10'd556;
					  10'b1000111011: reg_q <= 10'd557;
					  10'b1000111100: reg_q <= 10'd558;
					  10'b1000111101: reg_q <= 10'd559;
					  10'b1000111110: reg_q <= 10'd560;
					  10'b1000111111: reg_q <= 10'd561;
					  10'b1001000000: reg_q <= 10'd562;
					  10'b1001000001: reg_q <= 10'd563;
					  10'b1001000010: reg_q <= 10'd564;
					  10'b1001000011: reg_q <= 10'd565;
					  10'b1001000100: reg_q <= 10'd566;
					  10'b1001000101: reg_q <= 10'd567;
					  10'b1001000110: reg_q <= 10'd568;
					  10'b1001000111: reg_q <= 10'd569;
					  10'b1001001000: reg_q <= 10'd570;
					  10'b1001001001: reg_q <= 10'd571;
					  10'b1001001010: reg_q <= 10'd572;
					  10'b1001001011: reg_q <= 10'd573;
					  10'b1001001100: reg_q <= 10'd574;
					  10'b1001001101: reg_q <= 10'd575;
					  10'b1001001110: reg_q <= 10'd576;
					  10'b1001001111: reg_q <= 10'd577;
					  10'b1001010000: reg_q <= 10'd578;
					  10'b1001010001: reg_q <= 10'd579;
					  10'b1001010010: reg_q <= 10'd580;
					  10'b1001010011: reg_q <= 10'd581;
					  10'b1001010100: reg_q <= 10'd582;
					  10'b1001010101: reg_q <= 10'd583;
					  10'b1001010110: reg_q <= 10'd583;
					  10'b1001010111: reg_q <= 10'd584;
					  10'b1001011000: reg_q <= 10'd585;
					  10'b1001011001: reg_q <= 10'd586;
					  10'b1001011010: reg_q <= 10'd587;
					  10'b1001011011: reg_q <= 10'd588;
					  10'b1001011100: reg_q <= 10'd589;
					  10'b1001011101: reg_q <= 10'd590;
					  10'b1001011110: reg_q <= 10'd591;
					  10'b1001011111: reg_q <= 10'd592;
					  10'b1001100000: reg_q <= 10'd593;
					  10'b1001100001: reg_q <= 10'd594;
					  10'b1001100010: reg_q <= 10'd595;
					  10'b1001100011: reg_q <= 10'd596;
					  10'b1001100100: reg_q <= 10'd597;
					  10'b1001100101: reg_q <= 10'd598;
					  10'b1001100110: reg_q <= 10'd599;
					  10'b1001100111: reg_q <= 10'd600;
					  10'b1001101000: reg_q <= 10'd601;
					  10'b1001101001: reg_q <= 10'd602;
					  10'b1001101010: reg_q <= 10'd603;
					  10'b1001101011: reg_q <= 10'd604;
					  10'b1001101100: reg_q <= 10'd605;
					  10'b1001101101: reg_q <= 10'd606;
					  10'b1001101110: reg_q <= 10'd607;
					  10'b1001101111: reg_q <= 10'd608;
					  10'b1001110000: reg_q <= 10'd609;
					  10'b1001110001: reg_q <= 10'd610;
					  10'b1001110010: reg_q <= 10'd611;
					  10'b1001110011: reg_q <= 10'd612;
					  10'b1001110100: reg_q <= 10'd613;
					  10'b1001110101: reg_q <= 10'd614;
					  10'b1001110110: reg_q <= 10'd615;
					  10'b1001110111: reg_q <= 10'd616;
					  10'b1001111000: reg_q <= 10'd617;
					  10'b1001111001: reg_q <= 10'd618;
					  10'b1001111010: reg_q <= 10'd619;
					  10'b1001111011: reg_q <= 10'd620;
					  10'b1001111100: reg_q <= 10'd621;
					  10'b1001111101: reg_q <= 10'd622;
					  10'b1001111110: reg_q <= 10'd623;
					  10'b1001111111: reg_q <= 10'd624;
					  10'b1010000000: reg_q <= 10'd625;
					  10'b1010000001: reg_q <= 10'd625;
					  10'b1010000010: reg_q <= 10'd626;
					  10'b1010000011: reg_q <= 10'd627;
					  10'b1010000100: reg_q <= 10'd628;
					  10'b1010000101: reg_q <= 10'd629;
					  10'b1010000110: reg_q <= 10'd630;
					  10'b1010000111: reg_q <= 10'd631;
					  10'b1010001000: reg_q <= 10'd632;
					  10'b1010001001: reg_q <= 10'd633;
					  10'b1010001010: reg_q <= 10'd634;
					  10'b1010001011: reg_q <= 10'd635;
					  10'b1010001100: reg_q <= 10'd636;
					  10'b1010001101: reg_q <= 10'd637;
					  10'b1010001110: reg_q <= 10'd638;
					  10'b1010001111: reg_q <= 10'd639;
					  10'b1010010000: reg_q <= 10'd640;
					  10'b1010010001: reg_q <= 10'd641;
					  10'b1010010010: reg_q <= 10'd642;
					  10'b1010010011: reg_q <= 10'd643;
					  10'b1010010100: reg_q <= 10'd644;
					  10'b1010010101: reg_q <= 10'd645;
					  10'b1010010110: reg_q <= 10'd646;
					  10'b1010010111: reg_q <= 10'd647;
					  10'b1010011000: reg_q <= 10'd648;
					  10'b1010011001: reg_q <= 10'd649;
					  10'b1010011010: reg_q <= 10'd650;
					  10'b1010011011: reg_q <= 10'd651;
					  10'b1010011100: reg_q <= 10'd652;
					  10'b1010011101: reg_q <= 10'd653;
					  10'b1010011110: reg_q <= 10'd654;
					  10'b1010011111: reg_q <= 10'd655;
					  10'b1010100000: reg_q <= 10'd656;
					  10'b1010100001: reg_q <= 10'd657;
					  10'b1010100010: reg_q <= 10'd658;
					  10'b1010100011: reg_q <= 10'd659;
					  10'b1010100100: reg_q <= 10'd660;
					  10'b1010100101: reg_q <= 10'd661;
					  10'b1010100110: reg_q <= 10'd662;
					  10'b1010100111: reg_q <= 10'd663;
					  10'b1010101000: reg_q <= 10'd664;
					  10'b1010101001: reg_q <= 10'd665;
					  10'b1010101010: reg_q <= 10'd666;
					  10'b1010101011: reg_q <= 10'd666;
					  10'b1010101100: reg_q <= 10'd667;
					  10'b1010101101: reg_q <= 10'd668;
					  10'b1010101110: reg_q <= 10'd669;
					  10'b1010101111: reg_q <= 10'd670;
					  10'b1010110000: reg_q <= 10'd671;
					  10'b1010110001: reg_q <= 10'd672;
					  10'b1010110010: reg_q <= 10'd673;
					  10'b1010110011: reg_q <= 10'd674;
					  10'b1010110100: reg_q <= 10'd675;
					  10'b1010110101: reg_q <= 10'd676;
					  10'b1010110110: reg_q <= 10'd677;
					  10'b1010110111: reg_q <= 10'd678;
					  10'b1010111000: reg_q <= 10'd679;
					  10'b1010111001: reg_q <= 10'd680;
					  10'b1010111010: reg_q <= 10'd681;
					  10'b1010111011: reg_q <= 10'd682;
					  10'b1010111100: reg_q <= 10'd683;
					  10'b1010111101: reg_q <= 10'd684;
					  10'b1010111110: reg_q <= 10'd685;
					  10'b1010111111: reg_q <= 10'd686;
					  10'b1011000000: reg_q <= 10'd687;
					  10'b1011000001: reg_q <= 10'd688;
					  10'b1011000010: reg_q <= 10'd689;
					  10'b1011000011: reg_q <= 10'd690;
					  10'b1011000100: reg_q <= 10'd691;
					  10'b1011000101: reg_q <= 10'd692;
					  10'b1011000110: reg_q <= 10'd693;
					  10'b1011000111: reg_q <= 10'd694;
					  10'b1011001000: reg_q <= 10'd695;
					  10'b1011001001: reg_q <= 10'd696;
					  10'b1011001010: reg_q <= 10'd697;
					  10'b1011001011: reg_q <= 10'd698;
					  10'b1011001100: reg_q <= 10'd699;
					  10'b1011001101: reg_q <= 10'd700;
					  10'b1011001110: reg_q <= 10'd701;
					  10'b1011001111: reg_q <= 10'd702;
					  10'b1011010000: reg_q <= 10'd703;
					  10'b1011010001: reg_q <= 10'd704;
					  10'b1011010010: reg_q <= 10'd705;
					  10'b1011010011: reg_q <= 10'd706;
					  10'b1011010100: reg_q <= 10'd707;
					  10'b1011010101: reg_q <= 10'd708;
					  10'b1011010110: reg_q <= 10'd708;
					  10'b1011010111: reg_q <= 10'd709;
					  10'b1011011000: reg_q <= 10'd710;
					  10'b1011011001: reg_q <= 10'd711;
					  10'b1011011010: reg_q <= 10'd712;
					  10'b1011011011: reg_q <= 10'd713;
					  10'b1011011100: reg_q <= 10'd714;
					  10'b1011011101: reg_q <= 10'd715;
					  10'b1011011110: reg_q <= 10'd716;
					  10'b1011011111: reg_q <= 10'd717;
					  10'b1011100000: reg_q <= 10'd718;
					  10'b1011100001: reg_q <= 10'd719;
					  10'b1011100010: reg_q <= 10'd720;
					  10'b1011100011: reg_q <= 10'd721;
					  10'b1011100100: reg_q <= 10'd722;
					  10'b1011100101: reg_q <= 10'd723;
					  10'b1011100110: reg_q <= 10'd724;
					  10'b1011100111: reg_q <= 10'd725;
					  10'b1011101000: reg_q <= 10'd726;
					  10'b1011101001: reg_q <= 10'd727;
					  10'b1011101010: reg_q <= 10'd728;
					  10'b1011101011: reg_q <= 10'd729;
					  10'b1011101100: reg_q <= 10'd730;
					  10'b1011101101: reg_q <= 10'd731;
					  10'b1011101110: reg_q <= 10'd732;
					  10'b1011101111: reg_q <= 10'd733;
					  10'b1011110000: reg_q <= 10'd734;
					  10'b1011110001: reg_q <= 10'd735;
					  10'b1011110010: reg_q <= 10'd736;
					  10'b1011110011: reg_q <= 10'd737;
					  10'b1011110100: reg_q <= 10'd738;
					  10'b1011110101: reg_q <= 10'd739;
					  10'b1011110110: reg_q <= 10'd740;
					  10'b1011110111: reg_q <= 10'd741;
					  10'b1011111000: reg_q <= 10'd742;
					  10'b1011111001: reg_q <= 10'd743;
					  10'b1011111010: reg_q <= 10'd744;
					  10'b1011111011: reg_q <= 10'd745;
					  10'b1011111100: reg_q <= 10'd746;
					  10'b1011111101: reg_q <= 10'd747;
					  10'b1011111110: reg_q <= 10'd748;
					  10'b1011111111: reg_q <= 10'd749;
					  10'b1100000000: reg_q <= 10'd750;
					  10'b1100000001: reg_q <= 10'd750;
					  10'b1100000010: reg_q <= 10'd751;
					  10'b1100000011: reg_q <= 10'd752;
					  10'b1100000100: reg_q <= 10'd753;
					  10'b1100000101: reg_q <= 10'd754;
					  10'b1100000110: reg_q <= 10'd755;
					  10'b1100000111: reg_q <= 10'd756;
					  10'b1100001000: reg_q <= 10'd757;
					  10'b1100001001: reg_q <= 10'd758;
					  10'b1100001010: reg_q <= 10'd759;
					  10'b1100001011: reg_q <= 10'd760;
					  10'b1100001100: reg_q <= 10'd761;
					  10'b1100001101: reg_q <= 10'd762;
					  10'b1100001110: reg_q <= 10'd763;
					  10'b1100001111: reg_q <= 10'd764;
					  10'b1100010000: reg_q <= 10'd765;
					  10'b1100010001: reg_q <= 10'd766;
					  10'b1100010010: reg_q <= 10'd767;
					  10'b1100010011: reg_q <= 10'd768;
					  10'b1100010100: reg_q <= 10'd769;
					  10'b1100010101: reg_q <= 10'd770;
					  10'b1100010110: reg_q <= 10'd771;
					  10'b1100010111: reg_q <= 10'd772;
					  10'b1100011000: reg_q <= 10'd773;
					  10'b1100011001: reg_q <= 10'd774;
					  10'b1100011010: reg_q <= 10'd775;
					  10'b1100011011: reg_q <= 10'd776;
					  10'b1100011100: reg_q <= 10'd777;
					  10'b1100011101: reg_q <= 10'd778;
					  10'b1100011110: reg_q <= 10'd779;
					  10'b1100011111: reg_q <= 10'd780;
					  10'b1100100000: reg_q <= 10'd781;
					  10'b1100100001: reg_q <= 10'd782;
					  10'b1100100010: reg_q <= 10'd783;
					  10'b1100100011: reg_q <= 10'd784;
					  10'b1100100100: reg_q <= 10'd785;
					  10'b1100100101: reg_q <= 10'd786;
					  10'b1100100110: reg_q <= 10'd787;
					  10'b1100100111: reg_q <= 10'd788;
					  10'b1100101000: reg_q <= 10'd789;
					  10'b1100101001: reg_q <= 10'd790;
					  10'b1100101010: reg_q <= 10'd791;
					  10'b1100101011: reg_q <= 10'd791;
					  10'b1100101100: reg_q <= 10'd792;
					  10'b1100101101: reg_q <= 10'd793;
					  10'b1100101110: reg_q <= 10'd794;
					  10'b1100101111: reg_q <= 10'd795;
					  10'b1100110000: reg_q <= 10'd796;
					  10'b1100110001: reg_q <= 10'd797;
					  10'b1100110010: reg_q <= 10'd798;
					  10'b1100110011: reg_q <= 10'd799;
					  10'b1100110100: reg_q <= 10'd800;
					  10'b1100110101: reg_q <= 10'd801;
					  10'b1100110110: reg_q <= 10'd802;
					  10'b1100110111: reg_q <= 10'd803;
					  10'b1100111000: reg_q <= 10'd804;
					  10'b1100111001: reg_q <= 10'd805;
					  10'b1100111010: reg_q <= 10'd806;
					  10'b1100111011: reg_q <= 10'd807;
					  10'b1100111100: reg_q <= 10'd808;
					  10'b1100111101: reg_q <= 10'd809;
					  10'b1100111110: reg_q <= 10'd810;
					  10'b1100111111: reg_q <= 10'd811;
					  10'b1101000000: reg_q <= 10'd812;
					  10'b1101000001: reg_q <= 10'd813;
					  10'b1101000010: reg_q <= 10'd814;
					  10'b1101000011: reg_q <= 10'd815;
					  10'b1101000100: reg_q <= 10'd816;
					  10'b1101000101: reg_q <= 10'd817;
					  10'b1101000110: reg_q <= 10'd818;
					  10'b1101000111: reg_q <= 10'd819;
					  10'b1101001000: reg_q <= 10'd820;
					  10'b1101001001: reg_q <= 10'd821;
					  10'b1101001010: reg_q <= 10'd822;
					  10'b1101001011: reg_q <= 10'd823;
					  10'b1101001100: reg_q <= 10'd824;
					  10'b1101001101: reg_q <= 10'd825;
					  10'b1101001110: reg_q <= 10'd826;
					  10'b1101001111: reg_q <= 10'd827;
					  10'b1101010000: reg_q <= 10'd828;
					  10'b1101010001: reg_q <= 10'd829;
					  10'b1101010010: reg_q <= 10'd830;
					  10'b1101010011: reg_q <= 10'd831;
					  10'b1101010100: reg_q <= 10'd832;
					  10'b1101010101: reg_q <= 10'd833;
					  10'b1101010110: reg_q <= 10'd833;
					  10'b1101010111: reg_q <= 10'd834;
					  10'b1101011000: reg_q <= 10'd835;
					  10'b1101011001: reg_q <= 10'd836;
					  10'b1101011010: reg_q <= 10'd837;
					  10'b1101011011: reg_q <= 10'd838;
					  10'b1101011100: reg_q <= 10'd839;
					  10'b1101011101: reg_q <= 10'd840;
					  10'b1101011110: reg_q <= 10'd841;
					  10'b1101011111: reg_q <= 10'd842;
					  10'b1101100000: reg_q <= 10'd843;
					  10'b1101100001: reg_q <= 10'd844;
					  10'b1101100010: reg_q <= 10'd845;
					  10'b1101100011: reg_q <= 10'd846;
					  10'b1101100100: reg_q <= 10'd847;
					  10'b1101100101: reg_q <= 10'd848;
					  10'b1101100110: reg_q <= 10'd849;
					  10'b1101100111: reg_q <= 10'd850;
					  10'b1101101000: reg_q <= 10'd851;
					  10'b1101101001: reg_q <= 10'd852;
					  10'b1101101010: reg_q <= 10'd853;
					  10'b1101101011: reg_q <= 10'd854;
					  10'b1101101100: reg_q <= 10'd855;
					  10'b1101101101: reg_q <= 10'd856;
					  10'b1101101110: reg_q <= 10'd857;
					  10'b1101101111: reg_q <= 10'd858;
					  10'b1101110000: reg_q <= 10'd859;
					  10'b1101110001: reg_q <= 10'd860;
					  10'b1101110010: reg_q <= 10'd861;
					  10'b1101110011: reg_q <= 10'd862;
					  10'b1101110100: reg_q <= 10'd863;
					  10'b1101110101: reg_q <= 10'd864;
					  10'b1101110110: reg_q <= 10'd865;
					  10'b1101110111: reg_q <= 10'd866;
					  10'b1101111000: reg_q <= 10'd867;
					  10'b1101111001: reg_q <= 10'd868;
					  10'b1101111010: reg_q <= 10'd869;
					  10'b1101111011: reg_q <= 10'd870;
					  10'b1101111100: reg_q <= 10'd871;
					  10'b1101111101: reg_q <= 10'd872;
					  10'b1101111110: reg_q <= 10'd873;
					  10'b1101111111: reg_q <= 10'd874;
					  10'b1110000000: reg_q <= 10'd875;
					  10'b1110000001: reg_q <= 10'd875;
					  10'b1110000010: reg_q <= 10'd876;
					  10'b1110000011: reg_q <= 10'd877;
					  10'b1110000100: reg_q <= 10'd878;
					  10'b1110000101: reg_q <= 10'd879;
					  10'b1110000110: reg_q <= 10'd880;
					  10'b1110000111: reg_q <= 10'd881;
					  10'b1110001000: reg_q <= 10'd882;
					  10'b1110001001: reg_q <= 10'd883;
					  10'b1110001010: reg_q <= 10'd884;
					  10'b1110001011: reg_q <= 10'd885;
					  10'b1110001100: reg_q <= 10'd886;
					  10'b1110001101: reg_q <= 10'd887;
					  10'b1110001110: reg_q <= 10'd888;
					  10'b1110001111: reg_q <= 10'd889;
					  10'b1110010000: reg_q <= 10'd890;
					  10'b1110010001: reg_q <= 10'd891;
					  10'b1110010010: reg_q <= 10'd892;
					  10'b1110010011: reg_q <= 10'd893;
					  10'b1110010100: reg_q <= 10'd894;
					  10'b1110010101: reg_q <= 10'd895;
					  10'b1110010110: reg_q <= 10'd896;
					  10'b1110010111: reg_q <= 10'd897;
					  10'b1110011000: reg_q <= 10'd898;
					  10'b1110011001: reg_q <= 10'd899;
					  10'b1110011010: reg_q <= 10'd900;
					  10'b1110011011: reg_q <= 10'd901;
					  10'b1110011100: reg_q <= 10'd902;
					  10'b1110011101: reg_q <= 10'd903;
					  10'b1110011110: reg_q <= 10'd904;
					  10'b1110011111: reg_q <= 10'd905;
					  10'b1110100000: reg_q <= 10'd906;
					  10'b1110100001: reg_q <= 10'd907;
					  10'b1110100010: reg_q <= 10'd908;
					  10'b1110100011: reg_q <= 10'd909;
					  10'b1110100100: reg_q <= 10'd910;
					  10'b1110100101: reg_q <= 10'd911;
					  10'b1110100110: reg_q <= 10'd912;
					  10'b1110100111: reg_q <= 10'd913;
					  10'b1110101000: reg_q <= 10'd914;
					  10'b1110101001: reg_q <= 10'd915;
					  10'b1110101010: reg_q <= 10'd916;
					  10'b1110101011: reg_q <= 10'd916;
					  10'b1110101100: reg_q <= 10'd917;
					  10'b1110101101: reg_q <= 10'd918;
					  10'b1110101110: reg_q <= 10'd919;
					  10'b1110101111: reg_q <= 10'd920;
					  10'b1110110000: reg_q <= 10'd921;
					  10'b1110110001: reg_q <= 10'd922;
					  10'b1110110010: reg_q <= 10'd923;
					  10'b1110110011: reg_q <= 10'd924;
					  10'b1110110100: reg_q <= 10'd925;
					  10'b1110110101: reg_q <= 10'd926;
					  10'b1110110110: reg_q <= 10'd927;
					  10'b1110110111: reg_q <= 10'd928;
					  10'b1110111000: reg_q <= 10'd929;
					  10'b1110111001: reg_q <= 10'd930;
					  10'b1110111010: reg_q <= 10'd931;
					  10'b1110111011: reg_q <= 10'd932;
					  10'b1110111100: reg_q <= 10'd933;
					  10'b1110111101: reg_q <= 10'd934;
					  10'b1110111110: reg_q <= 10'd935;
					  10'b1110111111: reg_q <= 10'd936;
					  10'b1111000000: reg_q <= 10'd937;
					  10'b1111000001: reg_q <= 10'd938;
					  10'b1111000010: reg_q <= 10'd939;
					  10'b1111000011: reg_q <= 10'd940;
					  10'b1111000100: reg_q <= 10'd941;
					  10'b1111000101: reg_q <= 10'd942;
					  10'b1111000110: reg_q <= 10'd943;
					  10'b1111000111: reg_q <= 10'd944;
					  10'b1111001000: reg_q <= 10'd945;
					  10'b1111001001: reg_q <= 10'd946;
					  10'b1111001010: reg_q <= 10'd947;
					  10'b1111001011: reg_q <= 10'd948;
					  10'b1111001100: reg_q <= 10'd949;
					  10'b1111001101: reg_q <= 10'd950;
					  10'b1111001110: reg_q <= 10'd951;
					  10'b1111001111: reg_q <= 10'd952;
					  10'b1111010000: reg_q <= 10'd953;
					  10'b1111010001: reg_q <= 10'd954;
					  10'b1111010010: reg_q <= 10'd955;
					  10'b1111010011: reg_q <= 10'd956;
					  10'b1111010100: reg_q <= 10'd957;
					  10'b1111010101: reg_q <= 10'd958;
					  10'b1111010110: reg_q <= 10'd958;
					  10'b1111010111: reg_q <= 10'd959;
					  10'b1111011000: reg_q <= 10'd960;
					  10'b1111011001: reg_q <= 10'd961;
					  10'b1111011010: reg_q <= 10'd962;
					  10'b1111011011: reg_q <= 10'd963;
					  10'b1111011100: reg_q <= 10'd964;
					  10'b1111011101: reg_q <= 10'd965;
					  10'b1111011110: reg_q <= 10'd966;
					  10'b1111011111: reg_q <= 10'd967;
					  10'b1111100000: reg_q <= 10'd968;
					  10'b1111100001: reg_q <= 10'd969;
					  10'b1111100010: reg_q <= 10'd970;
					  10'b1111100011: reg_q <= 10'd971;
					  10'b1111100100: reg_q <= 10'd972;
					  10'b1111100101: reg_q <= 10'd973;
					  10'b1111100110: reg_q <= 10'd974;
					  10'b1111100111: reg_q <= 10'd975;
					  10'b1111101000: reg_q <= 10'd976;
					  10'b1111101001: reg_q <= 10'd977;
					  10'b1111101010: reg_q <= 10'd978;
					  10'b1111101011: reg_q <= 10'd979;
					  10'b1111101100: reg_q <= 10'd980;
					  10'b1111101101: reg_q <= 10'd981;
					  10'b1111101110: reg_q <= 10'd982;
					  10'b1111101111: reg_q <= 10'd983;
					  10'b1111110000: reg_q <= 10'd984;
					  10'b1111110001: reg_q <= 10'd985;
					  10'b1111110010: reg_q <= 10'd986;
					  10'b1111110011: reg_q <= 10'd987;
					  10'b1111110100: reg_q <= 10'd988;
					  10'b1111110101: reg_q <= 10'd989;
					  10'b1111110110: reg_q <= 10'd990;
					  10'b1111110111: reg_q <= 10'd991;
					  10'b1111111000: reg_q <= 10'd992;
					  10'b1111111001: reg_q <= 10'd993;
					  10'b1111111010: reg_q <= 10'd994;
					  10'b1111111011: reg_q <= 10'd995;
					  10'b1111111100: reg_q <= 10'd996;
					  10'b1111111101: reg_q <= 10'd997;
					  10'b1111111110: reg_q <= 10'd998;
					  10'b1111111111: reg_q <= 10'd999;
					  default: reg_q <= 10'd999;
					endcase
					state <= final ;	
					reg_en_conv <= 1'b1;
					x_reg[32:0] <= 33'b0;
					y_reg[32:0] <= 33'b0;
					end
				final : begin
					//z_reg[31:0] <= 32'b0;
					state <= (en) ? start : final ;
					reg_en_conv <= 1'b0;
					z_reg[31:0] <= (en) ? 32'b0: z_reg[31:0];
					end
			endcase
		end
	
	assign z_out[16:0] = {z_reg[31:25],reg_q} ;
	//assign z_out[31:0] = reg_aprx_z[31:0];
	
	wire  [32:0] x_sift_sign = { 33{x_reg[32]}} ;
	wire  [32:0] y_sift_sign = { 33{y_reg[32]}} ;
	wire  [32:0] x_sift = {x_sift_sign,x_reg} >> count ;
	wire  [32:0] y_sift = {y_sift_sign,y_reg} >> count ;	
	
	wire d_sign = y_reg[32];

	wire [31:0] unghi_it [0:31];
	assign	unghi_it[0] = `L_0 ;
	assign	unghi_it[1] = `L_1 ;
	assign	unghi_it[2] = `L_2 ;
	assign	unghi_it[3] = `L_3 ;
	assign	unghi_it[4] = `L_4 ;
	assign	unghi_it[5] = `L_5 ;
	assign	unghi_it[6] = `L_6 ;
	assign	unghi_it[7] = `L_7 ;
	assign	unghi_it[8] = `L_8 ;
	assign	unghi_it[9] = `L_9 ;
	assign	unghi_it[10] = `L_10 ;
	assign	unghi_it[11] = `L_11 ;
	assign	unghi_it[12] = `L_12 ;
	assign	unghi_it[13] = `L_13 ;
	assign	unghi_it[14] = `L_14 ;
	assign	unghi_it[15] = `L_15 ;
	assign	unghi_it[16] = `L_16 ;
	assign	unghi_it[17] = `L_17 ;
	assign	unghi_it[18] = `L_18 ;
	assign	unghi_it[19] = `L_19 ;
	assign	unghi_it[20] = `L_20 ;
	assign	unghi_it[21] = `L_21 ;
	assign	unghi_it[22] = `L_22 ;
	assign	unghi_it[23] = `L_23 ;
	assign	unghi_it[24] = `L_24 ;
	assign	unghi_it[25] = `L_25 ;
	assign	unghi_it[26] = `L_26 ;
	assign	unghi_it[27] = `L_27 ;
	assign	unghi_it[28] = `L_28 ;
	assign	unghi_it[29] = `L_29 ;
	assign	unghi_it[30] = `L_30 ;
	assign	unghi_it[31] = `L_31 ;
	
	wire [31:0] unghi = unghi_it[count] ;

endmodule

